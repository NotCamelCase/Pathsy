`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mfaJYDCVJ9tmCl1qOjTk0TJerc0+CZIKm9a/zNyIQ4axltn0gxS4ecX4Zo1Hni30YBnj26NHIuBB
AOWQWWIsIw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
fm/WgFN5BJ8I3UPgZJsI63Ae2cgM6RGTxS5FNhYU6XXXHkx0QJFyFRoU8CrUTLTBjuluj0orlDN7
b6tvmS/b+t2pz/hdtIzowwG7ASfmAm2Rz34QQjDzigPzCKTFoJ3AQFyFVp6APJAEpQMDshFJd1bU
o90A7irB+HRJlROZk6Y=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y9HW81s+G27R4EgUduReRfr2wwhFyWvK6LL9tlnP3yGocqrl4RiI4y+WWaJnw4C6dS3iiGHHmeJ7
BOLahMIyubxysrUfns7VGho/kNW6ikt7VXVZ5L5jmw9yuPTyIBFncC1xqSP7xNaS9k/ZAm5Lw55K
H315o/JmcCyyn5HSr1jVdFPIEuJ8RryEov/1F3wae5vQV+K2pdDVM4yhMeYiSV3rEXBJQCXsB+F9
U7k3P3lccYSLv8P26y2VMgzFU41xdKGkbGHUS4T0+mHvvMFy+vHD9LMvUteqPYdGOQNLjruKlAs2
AHopne8jFhsR31I7KARkwyENb8xzvOv8sBzGyA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
peROq/jTTnGKbWA0WQKdstqCMBnXCQ/l0MNC8U+wUBEgSuxXmaO6sZXlxNbYuvF5VqsLnRWixfy3
wh0htdw2Fg9D9Qk9/a80vu3uBTjVWr4lk8hrLkJnvtq2qtTfYk/OAyM32w2akdkxQ3wbWQ4k1AYN
qu5LIPFvpDfcjJlhCIKstIQm8wteJnd0cow/vDk3S4BJNKAzSiiXErh6GWgVub7ULXmltrFcrexW
PVXlGQKAGU8jNZpJxJZ1WZgcQMimYvj83x1+eJZE2cVzV8Ig8vWL+yju6Io7b1mfyOmpgUuApCtb
8AQsP5qESwP/N+mwguWx7J8Q08qdqM9x/QJkcg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o4FY5pOROZ9YI9RA5p0Ad3kE5yq0whzakHnr9rZ0OajyGLv1cnb96KSQ32j2VgDMft9OzYSZeWbt
PxyURKZ6s4QpIthjKZ5hkZ1dX7jaLHWszkXOn0aHalLo0oDQq0RSEei9uei7Mg0qW4DdwyOjJcD7
0tCjm+xUipiFJ626wm0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Iy13EbSeP18UOZBU/fyz/ghFg8ztq+t53D7w9iholnS1uDKpOjzlQvaeEBmYfRXs5NHQ14Pz3P9w
+hmZDs+uzw8iMA86Fp7fhnCuPzX8/LQRFToaDqPBMIYa6DRqM1d3Ld1ih9i/AYotsuhbtel9kyE1
dpbRQDO6rz2jrgw+W1kKiLC+9RfHxh4rhcUUxHELzdAKk4vXRmckDFXzxZPvws5ULUdbGjwbrHeL
iXS52T7AJBCxom553aM4p0xnK2cy1PSV3ogeM3U2F3Xun8eEJi4+tWr+CR1ygGtAA5TlCtAGBvlr
27svGBQX5xmja+iZxtHHExze4wnvgGrmhq7w3A==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
RVccda1v0fDhNCHInFVLDT++HfpYurc6dNEqM4kYp87QHa9Ne4fPEjHI+WvI4PAXowO6tW+feTX3
T/e5eJB6pzI04jJCjK6p/D781dDkkQoBKYIqxJbhmeoO2j84jr0MgmdQYY5cgbbaXIuN5kkFGQSz
Eo3VyGRYCmtfJlean9QS+gf87lkNNT4AKI2eG3SLkZXKRluUCldaUlqjtjKrif8h5fFZYb9yuwsq
fhunSKXAsc1KYi6QHcvOL/gbHo/Ilar3OtapsZn5TUt80BJZAKvR/SwXTTXVXymePYywgZdpaaY8
YYWh/hB3K51qvTWtnQTsDu2a/EjyqPwE0ZFcCA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ay7+KMhXAM+UC1xDUAyP7o3xWwNKph/1SVNJt0GsikZJSSnNHG4zsI8jvwLNjebEEu08CqdnL0r5
ysc20SPKfLvMpMvniIth+gIJXsmroMzwKRsuyL8YirXLf/GY8pGp7aLrsCvZjSURGqBV07M2Hnj1
d6antFfvhNW252Xw3orHYwuz/Lf2G6HLlPpILmo8finQj+mGy/O6EW+tu2HSFoOThajmRh6XgeYv
EtPqisdn40Bo5CRpA1oJxOuogvjjR7R4h19uU7NavRxTlXWAc9v2QpkQZeUvwwZSttxAMF+PjrSb
vwJLBacGapQwB5KVmd1Cw90/LnH5fHNhvEKDLA==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
qzOcFXO4O8zN9faGFsurU3eYSecabz3rm5c+LOHjNccH6vkSDJWFpMZsUESSlHQaqMhHRVfZdUS5
lGJ2RK9B+WPWUsy0ZigEqRrK8Qir/Anm/3u5fyCH1FzwryCyo7cm+I2k8+YF0SWIvHVzK8uvNd80
ibPe68fBwOAMylrWShcthBrq5gSqHohNeO8bcRihn+/rRxXxUIg3X5JdCLKA5xMLpnXPZtF81VxF
qBxhvKrrsPRjuNDEcRmff5TnFJffnST0IrV/Wrpgey+qfe34kPc/YnN7G4IcyDB0crCU3KGhkfiq
yoXrdivJtqDdYo5HjSra238d/I8AmW/W9cSGVg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 23056)
`protect data_block
hfxIkqXS785E+s5gvKSSuGp3S8ueb6sUPJtUeRRCyVAJp3mKzudFMO5ZR5JaLwcHOtS5Yguz2OAP
DYHUhpPFiMSDNcBAQufgVaoBJv8nmnd1tb60T2KS62Uo0ycJR7pRFXG4LamSTkQaDLHJp88jJwB+
w9paaTETVBhhoGlc99M1GLZHRL1ndHDGB19yRY00QhlDp5x4Dg5na86aOgYdciMklmwtSu8DPWrr
X904T3LQq4idxAvKWa7rQhdIA7BDYAc/zJaoCUIhKka+//5osG3mib97l31YSoRwOydYiTbI4Yzz
g7glK0SBXObcA7LT+t3iaBMKYwdPgTO6hVyV2FeYqoEruNV8pnK2koArcLwJKAdOUWXFLRMPAp+F
AfjHozIk+WTPTDQ8v4b2UO7Yw6LsnMfwnzOocUS+Tnlo16vgmpC97X8vADrwi0IezzAb/3NySgQU
pLrAgLouVLqMYhqZBUUuh/jfELCtYYBb0pTIOzpAFbPzh2UnWIpsEQJpQRFE80OCXG5FFOHDHJRd
Ju/3lTiTuWtIDwspYW7jh6aCqlHeHJMv3utbADi8RKSEHIf+s7UDzHQIzeUhKKP6gipI9vtx9nVA
vNcosU/3s5jJj5Xm2Togr5yWeMFT3sXqFt+B5Uci09Ut25CZrx5R42dGMwlYA06p0Op62WJ2nh8d
15hYKyTDafuP07FeKoWlwb0iDOHMIybSIFXpTFQV7gocyFF5srG8LhJV0zuWBDd3Wtv0C2LQuKRy
6LDMw3yDGyKqHDZghxKIJAIUMaXIwKXj3U8cb9JcDHfULHhC0QXOlkzY2AMnujw86icgl9d57Slg
+LuRVcWCgWQaphvFtPY2HTcx+nE5QCf6cQEpEVak58hDr7LmZe4o0pOrg5I8/t2rzIU3q00oppAs
9ZdF0exGWAQtG/7PiZh8INGZxGXU1PxRCm8hg65RUR8m2YPXey9bpxNitRS4khJmGonEmL7EqoAd
ZrMZec+GeItfj4HFMt7aKDUqrEaVzvfYvcmA9LPwX4aNahDJDedI6WdYKQ7SNHGegraXO6sfKVJt
ccYq7p7fMV6loSlgkrhElTpvuVwn4+6npgkhyECSiZdD9gEAEaW5FUgwY0/7hknngJ92bZS70RIS
9Av8llYCHuhAEDrJGuDHWpAf1oq6pvmYicl7+FY6SJFkPssocApH7O3YfTua83yhI8r9D4iwKfTH
2SqfM8rzzsTIwnXj66IhCtDhQVNMpmgW6Q/4v0PNcKZeEm63D/M1tyi4+UiAkwDJnisL76cePQEZ
pJbZ4/vG0yhPu39YqSbAK8+aDe0sTDfaOaYGpKAt1w6A7HK4xMSMZ/r66o/XM4yKRSZPXUobGO4S
1DTWQ6xScAxfXs69CcuYVnNPWXkUi6pyZGP6YtOZiwmJnmZh/IlkLwOYBr0utCA4pVmCrCtpeb4K
2E5E9IPaKvpjYHnrxGaraJWRZWcIUWmmIdTHVy42W/r6CzoAsDZkpwDYk8u5z1CjL+NWV1xr3pDv
GLAt/4R1zFqsuDlAWHDKBe5f62J+hMaFQKSLYl8B+AYl3c4G/Z9BoqwvAJUnXwZSP+pvhB9VB6EQ
zRQIOXw7T1sl6W0NDj4FP/agPdqNl8MSmJe0zPDA17+xqPBV9Ppqj3BDHMG3MRBAO/KOq4erddIq
IiQ54o+fwDQ1GemQdN7QtiYZnNMFOdIQrC4JaQ7QdaEem/upxT4f8ZaaobA6Kxvudq/3ugxbTtr8
seMPTzOvXDWH8ADJQBC5JXWnJyAz9aeixJCM8I2hm4OljJWx6yvYTQc4jXngZbUIoDeWQjoFcMoL
PRYWWx6018AXparYUr5X4+wyrk+CBqouhbP0wKZ24by7kWEeQJIkyf33Xfk5GgWo/E2izSGq6Rvd
jN0bU3BfTI4hwT7xk6RICUuqqiGj+WazBxdsK9oxg+Ud4He6nvcTL+yxzbEIChMlgks0BIAB1fxq
FAEJFk+ryyvVV1hcL4+RvQIkeVbSJFeKl5Xx0H++HXYa2B+UJcEeqv6GmXfu9nN265d2iBbbOuS1
0bilk23OeVMZJCMUTGiTwO05zSYZwveWh5m8gNbItd7P0fs3fiwUlhC9ISoZWG0BYT/ZiYHrp9d0
yhf96CKuXtsNqfh2wpI1IhhivRUsksaD/AKHDPrJ5CIjdLtQC850LlbzoovI1KgJNS1TgDRPvi36
TI2HTgRISWABJL06OALjyREgtsOzYqqbQDQo14QRrN23x6dw0FtKvLMFOZSJ0VYUV0scgI6MY/O1
2duKif4qXeSHwLAtlRQCs6bb1qXFjHpadZj+ZP5oB0qnFdAfINoZonlkONrWhuldsRUr7NSvCMWC
I07FhvDcwTBMtbg5AvddHfya5GOQc++Rja3GGvvCyecG80uUog2CjwSmn7z+POG0VvBTJ4jmp6mF
R0rSu+/Z8wY6LxBQcPC8CEMUKhmTRK+VQYImrZgvQdfv2ofQLL0Sal+nm7ueBxb+QiApn6QtCdac
OWDR63QSFo3Lg8RX6sWVdMRKqK7ZNxj6uUqmrmfrvz73FFRBv0o2/EQT6JM0pxkoYkSl/aoIrT2q
TobdfgU/dm/az64uf0aGLPemhe8fFTRrBfbyYlkahDl3EEbvq+Ww+DtdbbUIE7X5iHgNQnJkWqrd
sp4BG8plC1/jwDKfCuI/JKtAg+n+b31DFSFmaso9bzc93/qWAgXLNV/Ouol9+BD+FnoQOM51Yui5
/bFDpPPifj/Qz/NtgjBMydRs/1VAgkoUb956MenyMQ1J5BGQceRG01oOS1tfv0sXbHKGauKY0Uln
SupH+PhsFfrpUwZqefuGN/ER9nWoC264tcutvLUF5N8tq29OScxZwUBmmmo58CQ3MJ9sQJkoRl6Z
nA+qKsKaveGzlTdl0aCHDrGdq+FdeUjAxQ+DJPyKdiieDngng3NL5d54MnsT90XEsTNTEGBYdspU
OGYsVCC+YE0o+gZ/BddQoRTqoGLvVF6mZZ/JipJwPe/+ovS6MgYlxXqB8wE/NjuLCXFdY8ghJOoH
z3redx9RM1/0Ay4CF1S18A6z51HDBN9gCHwuulsueaIo3+IQicBkL0pyalhf94D1kgrrN0x8GK85
IbgWs3o+rp09rKJ8kSALwB8ue8fr8WcX22DREdiUlbPO1CyklU7OmY5vxAIrYUiImebuifhEsxy7
eiBqgAUj/r2Na3HhD4piTu6fQlRuDD1U/vHM611IV76NgMH59rkNbVi6Ie3XrQvVSXGyutFz47we
CO/yevh3sce8H6n57S+cWFDxGxPDkDQa4AarkWMCs1NgqH8umbXfHIRQWP0/CFz+6aZIOZAmkOF+
wJYht+yx6Di6XojZL3YU7bN4IsigaWMQ/REgU7/HuCaCc0Cix/+ltnPeaSSfOrfJB26Ngh4L6Kce
/3nt9P5PGjLr3Nd1tZSdbwpF4Ge0NH/GE/p9XncUWPhltvr6f6/bvjpVNBgdbY0gGcVBo7BE/rgF
M9GhrnYjfeHq0FNT/x+LVoCNY+sBEdfHfl+N3quqSjsxolbLQEyNouqQ/NkPx8U7j0O+CbUGDCms
7akqEXU3wF43mlTXzLbHt9LSrV7lFaX6Tw4YJcVkvCxSMNkrvb4Tnne6eHaaIH1lThyCvSmu3rpH
OUQ3KsG2VyqSf0GE0QlrIW9h7uPFJQcWyUC519mlWuxCNDCoxFxYRMV3OVcEQkNcU3Ajkg45oY56
y8LYpTVskfCFmITFNTzvgKXggpUfjC4gZgAmw6HJq7VgejxddD3OvHKPeDG+GBnJVXrJYHFMPlge
DB5M2UiqvuAOK+jj7ZfcnDrIBG59IVxl7RbCenXrmV0cNv9wt44hmbHL0pi8IY0doZgaX9Ti5QGH
ptOJP034YTHcTWt5TMeEZcEjKdC/3ZL7hcoWAG/kCNY3ZAqBCmJFzJ2LU2pvhdZ5s747aM5GBi0j
lze+k3PyMQ60sBdAoinGJYlq+4030w/wX/mqLKTUFQh1Kb4iBTR+YurtQ1uwNvdpattmW1IKgDWp
EbwEQ1os6BjM86ppYamT0kQ62kcdDSnmPRC7TXfkAAB7oOPDzPw20/ORcg46Yg+nRYEAUw3mTn3U
4b0Rq1+dcLP4JetJWU/2TwV2TBqzN1hU3GZa9q96bDdTUl2SgmVlZByM1AjkSPbd4IYyu4VEHiVM
zFQN+XKlA6hu926iUWEWzvZ7BBIK4lO3fCeq0dxVMuKOBvffzwxLpMo1WFXVFQvN1TayRs0WWhni
/bjwK3/viMnwzPDZHBMwSlqdZ6fhsiqm/QJmoFgeNXWuBtBSa/yn4oM+Vm0WDridEEkNHBdQQTCr
tCpw6PwLF+sZVYIW1oj5LFLRdjUrDfctnKzuYVf+/k2MLqRaaJ5pxxkHWImhevMd3Q76eKLpW7BS
/KjAv5bEW0ysQF3c4s3QM4aKjJixUcu31CUGazDgRumGBhrX6ZtNP2wvvQH3rhBS5x1fHy/oqcIM
WyMcQpk9xHKK9ezFhJS7dOoMqEu7BEjUZx2U9aizG6Dy3G1EeuEdOnX0m5i9u85XzFOtBDCFMaIV
yNg5R7YUG4AMWZR1OjE/20vue75AqIHdbRHFSeR2/JkFEn8cWa04+0aiijiIZGZBz1tfJZ88pYEO
P3IXyaobFmCo662mf32AUtBQxnKDKezLFHf5T7pHlGpn7dZ4rLe2DBH24Pz/v3iuclEAERzHNezz
l62HkFjYbIzX6gl2mgs0qOTpb44j0eZMkU8cC8yj+ngwHKH2rW3UdsFTtXnpI/Qs2ZQmhyw6QS9r
EptNDYXBfQqXXj0iV3V5XvPKVHsYBA05+idGNOY+u+79PsSv0qcdPVyGAbtXWikc8p8zcAVfj+Rn
SXYeg+lRbTPZg3uJRpTBUBi/5Enud/5Oxh/4IjnhSJNQCAxEYvtohEx0ECwJCw1dy4g6r9VyLQKs
zFzA4yDWyJ+3pm/7JsuY6tur+knjxJ7AF375fShRj4Oc46Hd/d/hmKnaWPtj+LUtLV9PbIxCyU7h
7TX93T7V+IYXMv2VSThrlPs3y6mLBT7pWL+f9ASeXm9K559zlFgrjOUU0qyuA+1u7LR+kOyy0NCG
ExIQxxmqzv24uJPpN/IZAEgm+dXe6JlTSTuPyJ2t2A7O/cM9AQUC/Xw1xjoWOt9WGMqdJKsnqCkc
TTo1NcSc5UIVnjWORyff7XF5YR7pChhIktfOTHsHO9sfJyvIxKO8/1IIKpWsx1PFIa5/EiQXwbCQ
SFHbFa2wiOWyNDAz3HQSxGfsZQcaH7F5j9tzpQgdnVDJrtGhBQCg8UNEUuTbkYp3j6Zr6GNIGeaP
52Yq4IjdmMaaqyIoqYl9CKL90FkK2kSRDVJMQRltlfeQwMK9rw49jdK4+ZYdy9uCmOXE8G8rZNfT
b/rMD3u9DRV2acvqlk1dcgAQMpOL4qGcQNCzHyd5JVpTFJk+mHr28hw3aJUIc+PYbnDk61I0si2m
Dl7YAXVQ0pFubFXig5i+YRj1l3uQHn3KcW23E6bap+sLEZoxjYPLmmCw62Z0db2oNgsbacnBn/Ql
/uGNQArX10YZgVrxkvlitatX556ZZhaZUiQ9KhUjJnqDwzzxZwKlehIZ2pWXPTfPzyayPgJCirgz
0+GGAB02gX3dutIiXd7Hy4GAuc/aUIpbeIRGLAkohjanSu8Em5m+Ta1/ZzT2xcbc/TtmuSK2NIUf
uF6wFZStlMjv+ny8DU7jB+0+B3SXGBtXtrSh0XdJcYPpggEiMWUD1WVyDwGKibweyX79CDgahKvd
nS5zsvzsHJlcZviw7LFUCNgY9g4XLs6MEBL/WQNYtKbDdt70uv7xL4GP6xmfddpM7Y6oQ62dMy6c
4+gPvHK6BpxophyPbcjwsoosrINgb6qywbyPvJsqeGvTt1AOp7snCB9ocm4eHAWnBHY+F5khJwT9
8x8UYIKxHFw9cL318AB9KU/8dXifXGanbj+ynqJPWnNfEhb5o5LudgjHf7yfBVGt4wum4vNjWpux
HkPYh7mVl6Jov4knCRfRVC00kXLAdrzH5q2q1g8oSB/STgfLbg7CIhj2PtIqcdyAuEj5tCr+j/lg
Ihr7UYfuOeVzMMgpFDWAvDDCO7W6lXWXNbM+bCD4TCWaLaCBDOKHbLaD5RTHSBS1mb6/bGJdJlcp
pzv4bP7ei9d4OEUtXkrvHJOaiPIIMTMiooyCRNXo+bQQOSOJGYpsZzv6gS6EIvwug8uxxJcPG4Yk
Q5rkrhtSV/JY56QQZ228UvUxNGG8WCrE/y/w87VzySF/Z3eaISKRfFuy+ymKzKTQYWouWkeuTXVl
jSqKVOJWr049V1J3H5GT9iOmGRb/+GL3pkO30+ENbMstzifWmht2qnXC7N/Y+oSfX9QL9EnMy+tb
r1yDDZD/QXfaaOHAhvP1qoBMJp6q/v4wRjW55wIHudP1zorCRKJp9bplBKHEDLexDYFTqGKoiVJp
FwGkmybH8IsGjo+hQYGRJv4abWJNzL9LJpGwAM8M3MDsrUZy1/Ai8G7U/KtYW1+6enL2RJj4uY35
en7BcCL07YyVdhbv5XnVCjVlmidEUZCjosEG5n3OJSlXUOBXW8LVoV0XufXwwP7r4oJMMylwt0gK
UaIODMg9qN9zNaKAKx5dr8u9DkDzfgCjmbAnIQ4gJpUU2IyheAU/gStVZVkeL36hxzfmZGc2/Mgl
lrSDUB+ezTUn1C5ogDF+sOy92qMC4XblBjwK5veU7qwNPwuZFC/BnSgc95lI0mdJqc1BzvfoWuLC
HFiP5Fkau+lJ36NFx6g1i2TvXQYxoQ1/tJZxsOA13egrG9ZTs2SG21rfydGrxAX3HSSfgvq8YdUi
rdlFUrz8rAARLfQJfk7AHPrkkPjNEKdvxZo7dYkUt62u8RYCQyq+yd4pcROwMgUMsww6BBm7wuEt
A/pS7fNqf2p5fia6P7bN68Vv9Wpcq0elA/LXV26gJo7EoZXmfNseQIMIcoXYZNtNQTcQaQeT5RXk
FupdNfDvckz85x8pcskj3xa1/+wDblrSelpQ4JBh9LvtSnS2s5CBi5SHd8CpK6qYCbbBSceKhG80
ka+vRKuVxiy1Raj5F9ClGgGHyjNvbLRuqvV7ljBef7P8SDoqC1GIrg/HME+gekxkntn3NEObvtE0
lICxcDS1lEdyJcU1EwzvCE+xm33fbZp18EJMD2pPwKbpF7mbBB9aLpb1L5tBikpFj48QPE65zoe1
HFtN9K5thjEZBVStUJC2tE1zBosbLsb8Dm0WY7ueo1dWTh0s99nL9TcE+ah3rOUUHNMWsTmDLozc
BRTdCUshUurEyUJO/QxstCiiv07KLvnCNVFFDEfn1RHLc2xS7r+jCgw/Cbch46ZBcZtux3cRi724
ptOzeFqbvt+vkabV5u2ZxoXygm1nW9oyWDDLJWKMkhwG2ADtLY6ZSFUO4+8f7+m0GXHTxuqWgso9
mB/th+BAIDO7zxcK3TDnVGKsrfmqCBVjIqvzKgJKwrYm7f+mw9T5IGNJTsDYJmOayBey6Uo8OVdc
AIdevWjfoIIkeMC58TJwSj0PhkhTnZdtvMAHuA2o+slji/2VAva9A8PotaPbJTEtjy1dHTySklVo
+2lYhcu9qpIStjdkyx5Yw/ISpSQxC0vws1wwjjXloBxWOjboTeiVt8DKeVpihtFegpzuleotz1px
NN7VDSk39RcKDfYf/8+B3qeJXDP3iyPUSilQ2lKRNgma7PLXxNfV861pbXBTUwR/W4P+YFpco57w
6YC7XnHofphxZBEKK6YnSufwMAVK7yTkHEGTof1AM+gDt1rzzzl/R+BiYbLf/tA0HGZ/4phrGVYD
8q1NfEdTUCLUZ7VJfWrgMGgVXGjJruLa6sI4sX0Tz7wDPw93nXZjljvecIbWq6l4DG72DL6q6wFG
Jc2hVPOGkusgDr3kQOYoF632HNa2BjpHJqS3Pl72Dvemjvyo2rIyu93wlh9m9/GtuJ1BXOwmb4nu
rwtO53UVPGu+x25Wa/XM2QXwapYFgN7UpTuJO3ZMabfgcwvkAA+NhSD/S6muhJFwXkMwx6j66966
Z8X6qttnD9bQRN6BBvruAuZMpwl1TRoS+Mx+ULrIFSwNbzZf5ZsjVF5rI/dzfveB/r7kHQj1nTpo
FDMM7sq2sS2wraVdAK+NiqC3AjcgX4hiAV8hrY6+UEEU+emtFlwA5hor+Sm960Y9VCWGHtAlahvy
dsZ2fUFWMF8eoe5m0yGuZFVQm/TpUY11WGHErHYAKpee6uF0tneukuzxd7L31jduQcGHTmZFvSkn
s57X8LSqL+hcSRzG9iMK9atnFqLSou3dp6zUyiOJl8IZkFBYDbCxVOG7xGi+39G3OUZXMmPXPfq/
BqMMn+15+NG92nn0IvCU2c9lgCdnNdbYZDtuupn10vvJ7mP/c+jcotNbMDWrQ8h+4r8kLy4K8tlO
CPaTXY+mPUTLYtDYP0xzIDP0Kb8NOPpsHNfoTizsF/4jdhlpC2ObQo40z+5+OtkEJ3z0n7JGa9MA
89ndlYzP0K6fT/PUC5GHMVb9oCH/stHMVB94DZjdHUOKex8ECHt+u7n5YE2ljEHW+7bFP7M/rfOy
CIo91S2kQovEj7MNVdMo+nJxhE7+xUPCLoZurrhxmH8gNNc5C5KqUPe5bHKZx/pi31LEE54Dftpm
YXJxKPLoRWBKPMtTCt/CVmGdUghdHsK2PotlI8vXpi9IifFd7GBP6o/28lQXUG0xti33tH416JJM
lLtglPUNunVCOTUhOWnRIwZebeR+2xW7WhjqtU1MhK3d8aoq6iQj8wEcsGvdAowG4JYhBuriyUvq
FuZQ+y4XMqTMk/bz2PzFeS3RKhCji4r2pYTGd5G+Nb5GqHXqlLjwLxoLr/RKdkjYYVoR7XviNM73
xsbQQE8/L6OpwfnKB+XdiDjJHUjjL8GoOOMHIWXuFq3n+QekrJAb/jGlmlBFW6aKxxg2sY+b2JT1
Dld03odbZac3BzM8W3QJyb/Cw3Ed9UHc9tUQ/WRcRGoPIRrQ6OHnncpXLxBZnxwS7HkIVx5Je90h
YoW9a79sK4cb5tZZGba2m2Je8v58httgteZTdLI8Z55oDEo/c6h80PzHMV/ZWMQqCFeV2JnIygeE
soIt+YrYmdyvoJKpQba5JZsF4DrgSSS/9tfmLk7chS/Jc6aFZgA2A9w7ZA0PB/QbvDqDVTvr46+3
B5uAT+mQ3MF9IZZXQhLksar1lwDHb92zvqi++sHgEr5zslyaimDwCvERobA3KULBNQV1O9glszqF
Q1j+dnrXJuGn+X1p05LqucA5RSnMao4SomfRVBSw00nyWuAq02/044fcQrtc15l9/rumHIk9/Hyv
9ypPB3Gd/cQjCq1gjvqBQuAL2xrF93KB+G4E08BjJDoT2MvIOMmtwgJlSUOeCxbhwu3izTK6IiVS
WUC4uIlQaxnOSdG6qokL8MhEiII4AMeQdUJfZd0+Vw9C+w7iQ4IJHl+YyCIDnfjrFYw2Hb9WqfIu
wnoKkRXbGrSlIN+qblDWJKqqvHDHVimqN8tARGOnH53hxc1/k4nI2AZsBtRtEG+vx0kicslH1GGM
aY1I9ql5R+DzUZCHmvhzGfXCgs0Ae+fpS3DDuh+vLAvSzrc+ifZ3YyH4vyOvQf7XPr/zTGIhjo2x
DElGh5pDNCYxQtfu+C7NgRfe+c4hYXLaTbGYZWViIeDybopz1VATExd9EkTdcTBnYGKiN6SSvwu2
lY/o/KRfLzxZSqZ4zfBCvYhIFdZY0JrxriOWEu5g3UWpvAfpYlrP9BiWtXVR+fookkZoEPPN+12z
3JyjhWvCskE+5SJUYezYAcqtel0ABoJJ76mtr7c7Jzt7asb6Rzl0AmOlXxLsn1ODEuDacOfhRU+m
zMRWPBLLCX9wW//THw3YYtVBsnJyqCbgpzz9UjQstlMfgLqAXq/awW1sKEwQ0nZtGee6P/entsZc
Ay9rvaO4l/9+KRNk05M3QwLl97o0eJHbv4r2K6UqMZ9G8fmDesDX/rkkg13eSzHZMYEZDI5Jx4Lh
iPqLT0RIxUXDM4DWL2L41XERARJuAEZcnkkR2O/cH9kzbOfjfUQ+1dYXPLi3dhUnYFALe6f2qVzP
aL3Lhzyivbx4DFU3F/Z2rT48yzfwvEIIF7iMJTAwcsMwA7tBiWJIP7xUaPATnPW+y4St8nSIUyLX
OG7bDvNPs8udU0NIaL5uZ2ep8dNQVJ1QjLD54MGladSXqEpTR8sS5u/vISpXp/QaErXtP9+y2jzo
qBfV+bWfMSuCqxEtcrqom+l6EkWAQVOlB9oIT8Q2lQWyOAz1qeQclgOCSQFLONw3GzOZO4noLbP1
QoSSDFFhNVtZCeq3WROjW86j8faLoS97EsWTaKWF/N9xhrPLbZqS4o0sDRSJCwGpA8GD2yaIeYMK
QMUaGqW37+WCmBjaw16AXor8fFDLevY1J4LMnVzASxuJoHo9BUIvayFWiFU9atEfB3uWKGaOLXs4
z+FGL4A4T2x7Fu1BYWB4kH8D/vwj7gzzCjY4jH/Qp/jZ2oYE5tamh91jJdq35qPhNM4K7AuJ4JoR
Llc0sU6n4SlGFkcgdrqQmVtl8zAvLHNRf9fK+v4yGSYZyeYMJeyvQOdCaNq7GCt0/jpldFp/7ozX
0ogHXuKwkMHWGDHVLcILxOlHpPiPIk8MF3L0D4GBTMdS7l+hdwP/E3hmOyYe42YU3lOyMpfGCJf1
vAryd93j+XE2zZ08jGOo/ikqsDZ/Gu57Sih7BNtr9GgAw/Pu+HGyyXLD5rfBAWdaip9WfvrOuwqP
+Rtab3rKnSt3xibUo0Yd1pcQO9SmV3BnW8UTpDPMFTobK063ARe7SI6/9Xbi4gKSN3ct3Ry0r8m1
kJ3YeYzhuau1YlrtGhzBKETE/3Qu8OKPSuDDw1jR2gKzr9yBx7ppbqDFltElElHS4Ykqe84In7Nj
Qf+0Atzbj3WTijBLOfY1ZU/7Gkj1siK8ad3FkIhAy6K96CdCukaXlJBp4icaHKSXKv9BrJKDyWZa
2SRJColCIspR61Hdm8XzmJfHuruQqI4asok4YIt0Q7GOaqB1LNjMFe7eXc+W4NDOElroziblRwpR
05CDLeYNWQWD9qAbn2Btq0nXmXRhxtID+Jxhw9MJTWVqo8tesGfc5zTcaoDUUh/w25+qp2AUmxNF
vnG3jMR7/4RxpIO4hhBVLqas80DGZk1OoQ4FdCHrIB+WVvp2gR8I85PwJHla1zFPYwE/1KgObAhV
tzveb95bMAeWEP8NkMTjR7w5EVE67wYSAeUdTEofzB/KQiAYxnBfBPqjcvREGrupPAoPRFUgCKSd
Y12rAKqgUOeBUDi/8M6XlRgznHbBosPCerrfwfQKviCH8dzu5fBW1qk/2rqkghJfoCiY6PDwDIDk
UR4WLQzHRYVCqv/xY7FRMG6j9WnYkdIDpVk7EEMk6GKh7jo0iLhmky7OfV5WlNWILvcuLPo6Pqx9
Zb33YhR3vH8t3Qe90rtkUupozPlpjNtoi8pPssvpFsrk79qnJxjc19kFlJm3+pIe0OlKipZKjUd1
Yv7r1pnobfYtznxx7H8vWePwHXCv44LNEFQHN7Bs1NxtyIIfEdSV730XoZJ1BxtOqsTSv+f+NRQ5
O/+t2Bg0q8xy9fy+TbLkUy9QK7YWwU1f8OWsxsJ9USW7dbbVRqYhXV0yP5dJptEWMHozAbc7MlEd
amljg5JTSCp0Icmkof5WjSPV6yImrU4woF6sWcPGJBOebFrb6xRpt45o3ewXs6CW2690tc3EmN9h
Dcf7DkZvYAqSJfcaA/L1p33SnPJPzeegimf2BaEUqjTXKsGCxL3a1GZU20f5kwktnxsRL+QoCWml
0rg5VTHhuyqmuJRZSerrkBo6wJ/fOwNaWlNfbqSdUTexN0Skn+FUiWwsqnp7x6mLA1nnWWJQCcW6
vNhwbN4GN1+oJBES11SCgRI8PLvS08JcNYT7+MjD9myTU4LRvGY00PGhJXcdBf8A/c6SM51JRPaY
lbvd70Kmkq7r+TYDgCkiiOB0goDheG0GBfLYfi3znpdptegl/SNjkGLXHbrqfrhvq0eCmDcLnT03
921+ogdTkb/F6Y7CA86IGBmzrNXXK9A9mXCR7eZ8SwUOkA0WVgs3aeFoWDARwh6PeirmSaoLi6u1
hyu5Wi4zNnhsBvQRWtJ1ZJ0fPJ4wt5C7vlRBVUF004K8AEvshxEzuQIDEAI/Ez2ipvSdYUFpik3S
mRyObCwBk5rh4gJoxXCQGsDsnsSLTIGhnUUSfnD4lWR5E7AcBAxQmbNVeM3sqt0xOSI81Pdrs2+D
IryexIwz5x0FzzuTS8MR6KarGWAyokZ0JKPLj3kuISSN7d21ZUM0nPc8roH1rMaYWkOj8Ay1EN+D
wjFJ8raQpqrS4uz5l2SpW6UikLHE5TAxs2OemgvUaPcECB3lRinrNjHsk+UzgYgxGU2vfnqr315q
pIh6kxZcmJpSuVqTT4yFY7Kwv/j0QBHZm4aLG9WaD49CkUFqBKfakl268DIAamAdWG2TEP3x3AjD
3tWElUOHMoKJEjOb7Mm18gQFDw4RszyL3fJvx6Ob2Dju/6iJQ1PJ2G6n2oDO45NXRZXk4S05Z6JY
IugjKU2MV5F4P+3q1FikEEA7lk+nN6bYNUdKLWqasWQo11uaVgV8USXiagMP1tOHqyxNsr533nI6
1gbSIJUex4Wfme7wSg3DFu51L2YS1mX/QU31VoPVEH+fVTBfHfTskVm3XnrRVd4OkZXLzVH93swV
QoCRls/KzTHMuekLcOVhbK6WUsF1+9+oLlwaih4woJLZDxNEVq/XkWLgnnSDmIewZzBsVHEgb1Q8
sP8HrhXulfX12AsOu33wD6Ky9TBP+cNKEzCdNA4cRHkOlcjwY03vY0o0hs6Y99O4Fq346UVHCp+C
SiS9O2wrBO3FF4gZjlf7V3X140yMPEG5vU37PsSDldio4yVAqZAlp0H1B6vhZwkwk85uwFa4zUaQ
x4FKPaXPkZoJlc1e6F4awMavqCneMH5kkhVFa7H+lrUpv62VzaP6ZaP/cDdiT7pjVACWKPCVkPws
IohWTxEWTYIrjZLvfhIWY9oHLs8Sc2Lz9kudPnDHKLYyN80sBcUZx70U2zvFgIOAvcjdWGXcHVcS
9v8hf3dfr387utrOb4N+8LJaQlKR+Cpio32CIo5JrNP2oigDH6gDfv89dnWZ2tNi2azCr5m1iZzb
zJUkzpiGwTg3lTWa9jMpyERkXWmXd7JGYKos8T7NQU6lxzdU6ySqH0HN9uUBEo7CypTbkLvCT9Un
GQ2Zdc7MC3gOuOmlPRd0Tn1wDzn45MSWbYWXzl/PTzWCqXMLx4RfR88LztNr7cDm30+nv11NL9uD
QN2+fNPmRcp3RIWF0WgwYKa+0TkaNY2BSjX0/q3Qzc/rX86rt75JDeD72m360+iePh90s3yXPFSE
bChQvxgVjPOSb3glN2DivZkbYBi+Uso+ax65FYF1Idr3gEkqLV5TozbYUiePg1YntIMmfglwVA5h
fFuyFWY09+zQxGDgl/fO/py8HwNUY77ZJ5RZT2BFdNnMewoPgNItKbFW+9Y452rkj5gaht2+tXHT
2gys952wOkS1IRMnURNkdDyeKm15pnQ4xe2MaOmleYNFKrz8cdBH82iCCVTiyiA7zOmCTqtfyhwq
wm86mRLuQo9j1BkK3clGZF89EfTnbyU7fmP8Yp73fJALiY/E8u+QbEWo0B3xW1dK3AyR4HE1xBbD
WfAc8JQpIMOMx0I1jmqJ+fvmn4YNW9wmBgaXdKsYWlQ7LoOZrhgvoVCob6navJNQCwGsrVQsBGNy
xm+TrerdHY/nF9w2h6KyVgwfNLrGC9xUYdHna15S1l9G0qseyOdh9VeReWX6ADEhbr/I1qp4JVaw
0SEmDgcVHin3wjVwKqQ7XHzAOBG8MvDAq2vVptRcYuAuY9flZHhA0sShFmi5qYmfXioST3Rm7Irb
zQcRlbNPmdzyRhJjzVcoY8/uUPZzHhm5xjJwzbGUKDZ91Vvj5b7t/NqKIJiSQpafB0WVQjd6KvmV
X/oy14t+of9t7DnH3uCdlHpCm48vpwzttXIjHFdTfZfoaCsrKHwA6ocGIIkIMEchbcRpnGWCJ2QA
G1cjZzfKHErX4kV9MYDkFs+3Aa1wOAIdJJoup+znGu+hO+8sYSrt1VzD/uAEHCWhKxmgWRGDekc3
1WifS6HYMtbBO7w8ZX8pwH+g0EiARUW9ellne8Thf75keshPoorKUd+5ph64jtVzHy5aadDLnVWX
PPODx6PTxFd8Umk9UQKq7WW+hDrvfZjwixP27N3Pcg1+jLrHS5wZxbTnmkkpCLfuCarR17jEM+8F
fvrlXTTA38ly1ljIRQbay09UAfjGtQVYXf2QE+jZOX5fZ2T+1ao8wVa3MwePzGvMJ6tNjw1TDDA8
gH67/WS290jO4k0RL8dTWwJEcdwBvGW3OAc7T85/V8c2qxHnbedZSoqaaw3WO5CeNNnnR47bZN5h
pBwzRQ4kk5rDS2/pNXfN9dDviHoD9e6TPphGlXBT0zhKCzxaau1wMOJN7bjhasEhwddiEdwub0TN
v942FMMB/6hKOt8l88iy/Z6s6aUrffJk+jKA8t1AdhkYwjZJsA/mZdymvV26ITOAVV6rAr7/Dwnm
1w2ACuga7/u6DLzeM6H7IcVZOWERTTrHrLlVPOh+AhQ+8/vSp1yyal76jqm/O3EYiAQpAcvchkUB
59uDtnzU2A3dDjFyEWX/zne2BSm2sfAyadiZFm67Uc7ndP2iDEXlaUun+PMTcm35mH042yPsZdSF
xN6WC+LJWUboAPAjmFj0g0L6oGEbdPE/Mcbp2uC94RzTOdyKzSvOqYXPG2IR4lTIpvIKVHk+Nx3j
/+8Hsi4FqzuNsaajkBVI1fLYQprsOaWlyFxgXn5kEekph0IRjT3Q8o/cEW/6YSUizlDFikjQ3V8p
zCaUbvgmINGswJI71ph8r+Wn9nxlYsDXj3/jW7cX1BqeTIFOPje97HKzimGzWCQAdexLkF+JgqCH
cUDqNLkzwYha0T2iHVUyOrcqJZki9CkpbCx8sni7vsBSX79owq+tqIxvql7rv33n6Ft31zEXG3Lr
hRsaZ0BZspMtw2P9sTxEV634qOj5qud7lmXluCrh1l3H0blkYUGrwmVWjeNbeT4cRxZbOG8L0+mS
ekvAeHrCDHIfsCS3sX7N20dKJU77ftR8P/SrHftyjrl77fWyfsLUsFg4DgS9nLz2l17r4iDuy22S
tXyGu7GiloX7myHlw5g0xDcEUpoYIDE72cQyqs4f/JySusgWWoCQdxfydhgdFPPxZgdax2d9MKzW
2PbG07Dv+3m6/i6imcwqrhRvaATIYPOesv9bbKu5v2NLAIUZTMs8TKOQe0gJSJcdKEc446RDuEoV
ZugZr55wcH7LvCmIH1UahMh4sc+mH0Q3X28WsV3/5PqtqdQJprQelZBXKrGgMKAL7rQCEsaQPhdG
xEWZCDyTDeoZObtQ+5X7MYUUHKEwQ81lkQzLzmiQ8NtsZ83XGjjm9My8Dr3chkbhmp7kIU9t1Bj7
Db4CFRcQdW1mf79rEXzFdbqjdeyenC06xLF2PVpMhomk21bTSd/K0INEvjeQBUDp29DUjY1t/9/9
TCN90d/LErzoKgdg5cOsBFmaCeLdDUVHuoqPlYcnF8wr0XYGoA+QW8yVUF0zkItX3L+9y5jSbBTN
vM6ePJT8rp10XPDvSA/S6KNdGnIdXfmwBSgVbwc3W4naaRu7xYvk17lR3n0snt9bOnf3zuF/H+Bj
a7bdFDxuWgnQOe4kJRD24ij7gioU43nw5y+VsMtdTabmR4hNYJ63yEpz4lVDIVBmxTPYBPs5bh3s
Uz+ZIWqS+uZ7M2dDDv/lyDTkrbznP8t1OlVmxfYQM7GVSydh7LVd7jSpVnMaMFMqVsek5vAQSoVN
eKLdTQOZqlIyQtMJSuXGSvlqjokcpkJeWwfPvoUwGhj0l48ybQdaqg7qGTch+6a3nMxipqG6e3k2
GCJ9/onqMF3oB6OXaAUXrfiRrO5jCdqI+MMyOF2JdnjNWalDU3OvJXBjmepeP4llq20Gopi+n0LO
FpErZC0ueK2k9KEKJ/xpKt21vPDIML2xrEGOK13RyAJ9wWc+0yKIKMtg4wmevPtuYqVHNDsdJI7z
bFCsCz/be7Qc+k4psxav1XLcvHzgqzwFHp3VnVdkz9uBFzkQehrNi9MP3p538Uib2JCSJLGggUkU
/7s7UGnKXXnUuq9znXYZzEiYFZ8V4QWvgfevfjfhcbv1DhY98NHkeTkOGY5JAmdok6gRXqyDWtWz
y54UqA7abC5/BKh680mkYLZwASb6xBNEX3Hedj+Sm9S51qhBvYxUtago8z9bgTzKJLU7vEtTLQlo
wytp5BYwFikrqR4N25U37K9pmfqJSPG42LZNgMgSk49ylH/wWZDtnWf8wShk03q1seNq6QlyGb/F
sTgNS86XR2XC13PpNP4vEfi+IhhxMdNWh4k2t83t5KloNRi8X1QqtzZ7OoZPgdrQRUQgr3x1WVJf
iD7BkU24zn0U11HEcBFWgYnwevvtpzXEjVIrFpvSjFzBSaSUEu5TRC1gIja6ot7GGAxSo16RXaY5
t41lWZ20PlSx1aRi3ajN7xAKsCAmFINpBY2jaNyjIWE5ujjKdcRTv9L1v99YwBf+nSaxaXCQ1xFN
YelOn+eRjfiTdkKgy4l7/QrpfjNUvi4zF1M7YSwRAMkamWqIs7mVfOGrILscPHivbpOIsrYg9f1J
YW33HbF5TV8daR/QOcLyT5AtsDgXO/3SR/YQ/wA61H6q1FE8U9tFrc2CuWnDHAnqHgFDrrDRBUVl
KM9R7y2ANq8M4cvFRhFnNXj4ELnnWhy6OXuMDsouR+xDqoI29/0W0SfnK35EUcRinTzjISCvtpL4
rQQbdxwSpJ9bx1UCpTSaKIzXzP76DQpntNAqEJ1zF5Rb0z8qvO4PZ0Ia0RACelSFU0Pwk/X333ho
cEfyNQhFbnCsWLAg4lXA2Rs7HVi1H2HuUxUlvdQH4IbKFBM/24KqJFSebvNfPNza6b5Zb4kXEytA
SDTy4T/VAyuoI0CMw9vjO83ZM19VpX0zfEwPbT4VYaci5TL4aBGYu1AhJvm5J/UkMqSkj728CjcK
ntiqzBezEgAZsl5dZdeFTahwjTROIqKl03G4HJ6x0cMW83CwsRPJXsyZXI2yJMqwo77t7VWdSK9L
K4Uk9pwMY3nUqRlJwP3e5GxhaiLuRtREpEFGbvfu37VFQXk9O8FK9QK1dFZNfU+nmOHAsmuAO3H/
PG5wbU2jnOiN5Cevsx5koRCVGP4cgjJFHz1jVMaVdxxGwD6YPj1Yz9wcFYikBMOG8cil5B03X/Vj
w3gk1XhlAkzpjeRx8xEbHZdiu7m1F61Ftk1+rB0LZAYYL0jjuAhoYNNDVm9/xaMQar/zoIt2l/WF
NMrm/xrELajdeJ38GGY4EFTALvh34yT+48iy0h4u/QajM9qoXBhKDvWddBMIe6LmUuvNginSlxRK
vWzescAMc54/tp4uze7WBv64GI+bIOWAOe/33f5Maekdw9irHnk8GWFVs1BRNF5ETG1AVBs5KEqz
IBdeJ2lxtQBtQKZ9QRJa06uYZTgBhiOl2EG6ADL2iyWQR5HIum5wVCT99a91mu5MMDAVWL4DplNZ
ChIjWPl2vdJ8hYLYGDLd4zFD78xdMvQb3U/GgO5s6++TKRp23OhutrEVdf9JzLVEsEiwtgakLQUZ
q7cNBW5QArK+USu+pNnOzRZ/VgohufmeojkdQqDSnYbHmUoNb0nBZU3L794AWRafe96eBGRFaOlz
Ckp4y1ao5BnMAtTtch/yPwueolzxevMxPi/MXKjR3gqontpPhtaJteR4UaGchs77pnRT8hPkepsJ
69PO26NthVHewS7pip3Njbm8SQg8BuJIjfuXpEj4603DgeOtGR9UzrHzWjt/ukDgUGqSuJmYcUAM
xH1NjksqTCdvFV7vf8H5PSaKXwDOu4vHDqcregTIOs1edDvUaCvcQWMxR6z8S6amSDnrpSANCL+a
wIO1GaSUwVDl80XpM+u7EkmXeVAQ8XbO9mamCvhvY6YXW5wQKKGC9qS5y5TYYQiD06zhLDvPKaqI
T4ttJQNH3CNCKLz1vKOTOm7hXFZFBKueRLtjrThWiL3rEK+Z+/YNxUa/njQZ2p2wUFm/TKxm2G9l
hBVmzKil67NzCZNC3JW2egSl67HqoRwaLj/LcjBUmsyB7mAqOSSZfIvfff+hEYrQOkl2mhNltlrb
td+9v2dvNfKBYYaMOc7iArIVLAG3NziiUy5+681GibVoTb9e/0qBW3VAxlnBeBeSBsIbGf4cbkeK
54TNAw5EvJlPmlm58F0W0KLr97NDUS0z9C3JAvFaMbZMw2lpKUjgGAT69wwiTOA9jUp/3xfxnUwg
bf6f5de2brX4dRMhnJOIF6/UqZSsucK08T0Isr2DcKDxOWrlD+MrQ2dhEVARcp5iHXNGcIUgTULP
1a6dmokm65EpnIsOQduYVC9CKfTTCjCo0lt5cfPlwhwnfp8RH5a7UEHoQWcScW60NhtB9MLP1Y+I
eHDBpRBp5bFXjpiV2sHmDObb8RD09BrsZ6H7ZFOUJw3FLm8VgJ7mMear0+WdcdwhR1zaYT+jeZkF
kpYqpAoBCMJ/0Unf8V2edcQDRZ+yBHcwvDFJjmBmpLZ8H7+KTK31wGh6ZvEZLCMi09OMF0WeMJYT
xalA5p2MgmEf3ERLyYfjmBVdjoR05ip/BgDjiAsgmhIXHg76/Zyw/jj/PoPwnbo6s3uRDWv/5+ac
EBkwa23xwu5LpEmBpaW2gT6uTMnL2cK1Sbi+KMWcKbcTNFaUnc7zgUoMfGsA/u7ixu2X0Tsmvm57
wdonWbqnbFxo6wZBc7P3306tZtpYVLPEfDdc0VRw/3fZOgkYDpndcUdXIPX9JVQHBtGQufd46Z1b
GrvLuLdo0wAxuCN5LRfKKVm87dIKPy0VjvElcUJOvIztTtr56dWcb5i4ALkKFnl3RCrn4ED66T6q
pPCrlqCW5E3ZvSDTvgS5v0HLg0yrrKKaMcScj21hqyUOjEScNOAluuaaiGPHdU8BCCeFYkHzEHHI
rvLAwdMKZGFmm3HOborH8NLuvazmL9pNYp5dFMOSpgqFQDHF9JG62BbTNPIXtJYY/b0v9T7zU/hn
3kVBj65sTbuz4gWSASBdRRk04SmDlyr2SEfGiFQqMRebsEQzyTSgTDpb4JuWZ/44J6HOfIrhoH0o
7LElmNPVkCYi3Mc4/43/KGkUqR6snLL4TKhSGUzJrDILrMg/ulMBZ6ymFVBSqK4heVSD6wl45XZ5
o1GAoB5xyQWqycrnq3fTYimFNmxYtCbTAzMWPv9jt4P5IlsVds7enzqVdo7zP+1GawQ+AKbokq9k
BCDlF1knEby7BtwzF2IDcctHL6EnlcYpJ7ICUU4j7Wdj/QBxMqf7rr2gxh0i/MI0SDdNUfRzA4yR
qXHBlAISA2hMT1yajmQUdyU4/vn0xAGs+bZPLTA+MALwQNlC4tqihW6jXfHpRtZYNOLXaQq6g804
oWHXLenb75BguzLHJL5ZRp7DQnZOeE/BOIyc0GuKK3XOgtd6CL9+a46EZc/O5UfFwD8kDwM7+4qj
ngxToHGv1ZPUurPMd/tewBpWa11c2yPlh7bQfeoQwHdDbv1xAmRqq66vibqjCy4XGPvPrQE3Plxk
SvMOdYakFxvtjuoJGicQckrp/6s4HBjy7eEoX/zuGObraA9yAdmNwn1w16M92H9YSP2detwe6Idu
KIe6wL2wY9jKWicRZ6ZCIcr8YkUIg4JUX0mYmH2xlAxQDc4pSYq4bfvBjXY++8YkKcDTWop5FClO
h46Li7j53U98SJktWKcwVD0fnbFvaLrK6zHUf0TfJCyZsSgUrHNoil1bDa4CD7nX26UdvsFlWEDc
9yLhNEmcCwkAIq3YlnogB0F8ReS5MijWUaaPbYjzSLguToNW3KmxBLocztsldJwBYaXsLlNtMQvs
60sLeTbIoCZ5FXQGCKN5kzNf79BchGwdd+3yjtdQ1Rr0XCiiR9WdgtZ5ye3m7WX+NiJkB/8gkKtL
/+++3cy5ksR28lADir3am6koeZ34cAE3FY+YH2Nqcbbw69KEjVfzDQZOMdMxF4Enh7Kzwql3Jthr
XENl4TIbcmi/QOSw/fDswL9Bb9viFLgIAx4pWjZ7NumOjN1RQIu3V5A3HF1xhZX1u3+JLhipJBC0
bpUL1dsspszxzlLLt+azrnzrggFTpTc2sDAzBjtXNGrW4c2kAFyQkWjePw2Uc8nsRYTlcy9TWgre
APqpg7BgF8IIjAUj8V++8vMswG/W7cskwrqMJnWoxJmgFDKf0w2IQtSLFkZVXhAFK4tiPbWFsedS
74deBxPu5KXEFFPI2yPQrNvK7gSdh035QrCZbJkYQko2vqJJDvbrQQxejQws0gwmOJEY+6rmzNpk
2J2HQHr07pPuXUKxyCskeiPcPjpa0dJCN98LUCpEJJ0uE8Q3/cyk2NkY3afcdG4I+0Fm6yJ2s5gl
jpXtebChiPCal8Uu7QOWEwRvc1uxJxzNuGH3FEck62Wew8TBS3PEXNm4ryTayL2F3Tejvh4U6ub5
wabjZrraYztQ0h8E5jD4RFvdqQ3qu0uV4naxE0lH3QWWHEaHEQnRwEMtZvdpX/C2FFFcSVCW5w+F
704LoeSP6L6+TgvedX4TNkOifCI2Z/LRAaDtfBEtzgFChdM8aQJhFF6zF+wM/PODVY2qlg9Alvd8
5Ac+Gr5MB0iRkyilBX844PYEzysQAZjdysIb6elLWZhgCuIq3MBXYL2emSQ4W3iDuJ8BN/djOw63
TH4u0m/JrTJQrA83SgEqqNDl8vG7PjgNpCbvA8qBrn7Chcum5E21jVD+UJbygXYG/knzpCct1g/z
uXsxYRm0BJYRl2ytOhsZZGtTcK6eEFZ4G3FNQ4gbTgiSN5IoAwbPSVgLUIgtEBX8hMuXWKV7aJqM
m/EdB1WfAmKkYBGgnrZE92iJu3/LzoTq08o95UyIpRLEfaF288t55GVL1vPx7pKIpmILM3uMpryt
0seqjlQeqngSkkKqixJ1YPZGf+iZ7Oi24XZPNcmiWPi/U683Ngv7oGqnc5gYqIUHQq7WwNyVO+Mj
8N1eahzaoj0gfw9mwvhB9SA5znsoyCLm3MjwYKioQTIuSUufYVfO5HlXAKymmdQQwbbTCUBmjKas
F6ylkHp7j379200uPGcIc0pi9mhdhnHSCMJqksEPfHQK0YJRy+tk/MJqf3SmayRD/eQZj2iIu+a3
uiMyi0k9ltLGVayx0/7yOID3Sc3dpJKVf2q7FVY/tMJavdzaiDeJreOhCYTuQ2SiEOfYLmcf2Atn
q5QgJiGeo5ixRCPf47YaoVIs7dsFZRs4HAi11IHx8fYcuuiurbX7KFOJiQBFuSe3AFzYR6eVuWd4
TDHjC/+KIy+Rz94qb1Hds4BMYBvyWUOxJtSI0r+IbPVEZfJbVqzUEl8KMRC2UzXfMOEFayX8MPqX
xNcSI1+tAK0SBNXgcTTjz6fEzYSvb/z6G4PyISpUxTNodUH5NguVGTVSgFBiFjI3FRxCHQKvnc8g
4I/E5RG5iBJXREawqSkybrNxqgA7Um0jC8p9rqmsZsZAga8ZeSx0KrtcTNqCpZgk5dArGLf+Htp1
poHYk7ccw6pseXelXw66HYh8/pFAlCWKTOKVmeXI5R+R22qyql/OBLaRq4JQoyBGCJnulyYnfFwk
rxZnlTtDIW8ufazxlhgRALUTYdbXJCLaf5AStaSiOnGgTZ2ODTmUXu3YQ+lwwml6K88au4S06Z/F
3+ZrbSRdC8XBduo8cM1p7Od2zdWLHeebzjWImi0zvtEQqRapV6HJj8wh20cAkpxe1ENmIEJl26og
o9HyWUwCXIr2RbmAIZVy1qduJteVSvzxZFSXgVGOeDjxHDvBjRTQd+0cKsezjPByrLro9broDOTE
l1bjfIzHXLPbsymSLXLDgcBJP633Y+eOk7cW1OiDlJg4Ztb31qjqV0QTx7UbSHfLN+Sy3DF9VYKh
7m+wS86+DfPpwjtMJkTw2UPcs6VmJGAAWtX7ABPxEGz9jBcV2nbmyF6FSS9hszNBw/8i5kxnsuqX
QG4576J8MJ3y6M4MTkiBoYS/D4VNLY0fwJN4oWnGzh/D1OnpfjvZDKf0jyhCB7ZQWfiTav2oSqH3
NQvo7a5RMRbH1fWsX6Xarksvgv5m88D1pvF8NKKkpXcE0PkMLjS0w6rr7Em+aYgwxxB9k+6d0JTC
XWu/eD74U+T9s5oUJbraXcSbddgNIWKzjTqpLsB4F0TAcGP51EZh265GmZ8WV+cDR+5GIoNl3pdD
LA97Sj/+xejCSrY08TIZUjOxeBLC/Pw3hnlxux3PA9lnk2sA7Sa+WUjVTYUd1kwiS1XpYoID51Tb
eXSUUFnw6z9/qePuKY9/Mh+ilB8/mOt5/U6CPLBZOvWGo+eK91aZJzsPIy32X+fxCYdx0xdqcGht
lZ+k5dfEy09VwOpLcdbbx78ury8Pvbcu4kD2a+F616OaOGzmr6Utloui2TBEug9o/cULMY+UbWDC
CHEez4lE0miPne6Rv/YQyH4sXGKdOiYq6PoMLk61tXlseV6l2YAKlblb1s1EQ8bUv1XSlbz2yERW
HNgBgJ/eUNrXmhR0DrLz+OHL6edvRfvE1h+4Kw2GHMF6tSg5l2SHXMcF5/+8nCTX//6biwCGdSPG
/ee2FcQyiu1wiaz0BkSrwU6nf4T61I8gTOyU7cVd7QBJ0Q9hfsqv5ag+wh7bDqqZBf4Dv7/2Hkq+
AujVzQqcxmND1f5k3JYVis+Ke0m8hhU7wlHjYo6C1V7TuVKEvGt6t6ux0EUDnxiDnN6yu3Hpv4HF
tkQztxPQ7nsdpnnLo5QzB/bX0fkSy9sRJCaEH6BvWc9+MTXXbKINviAEmNrZTGkyEqkh/VOrXveQ
PbTWLJ5zsMOrY/xelZPTzA2kZkCGWgejMG/Oyay7wgBUYwLb9wvC1PbAY/Zi/0GhdcWyi3S2yvKW
A+I0Sv7arwLPfeQzOMsAV4UYJF79UtN6WBkYhsETY05ka5ElX6BLkHKNQ4KrWvc3BTOaiPBsT68I
flhELAPBtmWAzZP1gp4T6aFvNvnUkSBoHBNU2WB7AS+EgJ8kbiBUg4RYfG06szQPuyBw+TEKP/VX
uom5H1dw1MWxt9tjxqnau7/3M3Ha3ij56kIseiYuEA/tjo5bXrVmulWWNntWSCUXAGwZVKAz0b0w
gEIR/f/hN9+0R+Ttvoy38UxNiuLp+l6N3jRC2YVBCiBXiPRkVduKdtjbCnczB5V6MZufvGwoO4GA
+nSDs7BBd+JOu6WRYhRoVfZcRHzNiyXrzjP4q10ceFYSruAm7/9sTn/cmS9CAKIfmErRqHg04+nS
rkSSE0chm+d/vPuIazDX51AfDUneuyYzalKEndnb6tUmbmsTwf5u5xc7AAph1oAGJOGZ4yzeAtjH
F4KkAvcyrUj8A8QVmgsxPbZ8Vp3PJet9A/iGIQIPCt/Cy3b5TguGUiSwyqgBTbTtVvvuiIfNHImn
d6SGLMlxTIC+gbAAuMYz4ZIN/cYfhToKO05MrLhhv7IBElYb8yl4YgjJoMGDiM/SeEEpvFXNissS
G82PidT+rRAexSAqt+/TFgTfyRZu78gwoh96ivDYBs3Pg6kSswjKVd7aKsBUzvYZVa4NPsnyhpYF
FZ/3t7YgaQTKiqse7cVuq1BRNoovdk8yV2ieDhcBrWoRG28J1xaCjzmcKzQpB2xngIwaP+ptnLp3
T46Q3euDieK3Uz2a1BE8wd5eE0QHcgly1alXifGeT12QUkIVLTyLCwjzzTaX2yZ+Cuvs1FTKIb+x
3nQU+26z7pN/uqNNWJWgLky+DbtObe6NtZvlA6zPq1d/pd4zkwy0vM1WM9gxnFdDU1RAMTBwWD5s
tEQ1yWFavT3G43BgCX1XkFCVn6Gdbb931kFuyJ3lRlyptezIS6qffakXTDwtNzPzlvRXI/MccJHY
JVuQ2rz5pGRs7Z+3bX2PzZJg8C2kWYIZD+Q9cS9GMcHShzZTn3dpQsBmOZgyrS7KA6MBDomd2BK0
u72foxY3DTlgaQX5yU/ROk2r2T5wrWem6hVa2Hj6NcQrF0JOdhpOIVxaWwU7OQW7xP608vt85ygc
cz9XLBXXKyDkQsvLSPqY8wkKyfzAJGYCh1BRr/+ylVDKGAOC8mSCdAK1+ixeU5UViKXTwgY7vK0t
DwtMgvZxYXSd7bI+z1p9nH/smyefXf0F90ylSmpMOA0JhbVxk48OmO/l7kdCLW2XRoaoI/jmGHvZ
xydolvsxzcr4lbOD8NSw/+1S3ujOuNhqO0d1hjA+pl12ud4vG2sGYseWq0kkTELZqnS20s5V9Y5W
iH4D379qQT9xQVZJ6AIYWorB7MKukKW1lNcJILoQFrBz07aFw2PfzTsHuVeNn0Hg1w2oVo53/o4F
bzuXfv2fW7WQsr8OI4zX2+k/boeJ+qB5AKxrdW8VNDpxNDlC6tfl3SQzrdaqWWl0Od3lpIQAnal0
8i/metbVIYvztM5vHFhdydtFGjOOr10SWRA5yq1qvub1wZh6M98nT6EkVYB+rUK0KE4co8AbaC1V
CtDrLTqzoGITZe1vV7C9gKYMNTat+txOtRMs4bRez608wsL/qy//WNpZgdQ9ilv8wKYzTsbzB4fI
ugLZXZH+G/QX0mt4V0YY2LTKNWJyNBWHnL2nLmV2hZx8xif2+/vUJXd75Ot3Avucvzjsy+bWFRZd
xGvFI97eBnMKCz7xd95FIdIK4o2s2yK+fdoFjTDSiK6UeJalP3Rfr9gxGjoTKXMr0kXDzDuPbgO0
Paj/GbtWutDUqLikYMcmI66IqNKvK02MNx3055LuptHr1H6O9WgZQw/4rmNW8aog7CJvBuoaoAbN
KRJ3saypfQfkb7jRRURDJQmTOYWKu8+kLBIKxqe3jRJAGg58g7pK+2Gsw86UOEkshYvaHXZW7mpn
fGECcodpfPdlBO8cr+Gz/jVmr3r3mz69uX+vIExpLJrubkc1SZ3mJUCeV4/yE33E0RY907O7Px8i
qIOLFwECSZtE5HbtyZN6LJDkSOBDkpI155iY4IxOICcuXfQMScXrSKdMq63EqGVxXpjAZmf1VSzC
zlhtZkJxAKL40RYDAw5paXz8sjUiQ6JF8jdMKLsjBigYt5SrGwM6eJf+iZuelvjnTTwdF1zaRIGw
Y6du33Lg3FKcv9EinIVStfHDdkIVyFz6YRqm5OeK6V0PrrcCkENmMTLfQDA1EY4qwFPpWzlu4dx9
Tv4anb0DZr4pM4sbu1T/JW1nZI0azCcIv3pxoJGDS2//lHsbERF5x7yrPyWJGRbt0I5XJU3FVpxW
iUrOG9SM5zxLL4yh6Lz9O2lScvfL5m1Hmhrpf8IXhqZMWSkKQbM5nSwG/OC6sBjURxh/xTsLt9tY
soIUsBEkf6s1hFdLeNzCu5Q0SyL3qyPZITvW3ai208XU3/VmQM+nezt56ie+8QrcW0xsSQi5kyWy
Jcj+SRIukCArzvD6NkMi0ZttCNsYnPUSgtMxmr6wkRhsSi7WEgbiS7fL39pKrwCVGYzRIFQbBKMa
WCUwHP0/emWmyiBWIAWY79sSuEJ55jYLA/HFGq5QcNBij+iKOAiLQRyyFRgdYxGWQbJzWDgPO4YE
c7+9wSziSnCAD1aqJ/r9mlryd1gdpcBzF/GJ9EVib6SU58z+x9W7O++5pTv6GNNStvM2go2VtBaS
1yqu2rcnMCC9CJonNlTdmF+3xGerI4giflpk057AAS4IJBrrEMbqEifIrKor+MuJej0WdAilToXQ
oO2JXf2zMjn7ViYC4lLq3PnwaIGHnqoqq4kz26rNlRYnb7SW9gKTGDcVBUdhU6XhOaTvLztd0PkF
jW5JXo/lzsP4nP4RBwBtMfWnJZ31Xum3kzshc2mkR81VJUTO19CJ64iLnFzbN1V2IUo9eSE2PTvX
FQsA/dBFtL3wXZBYaSVE0CHPphF5brDJZKKoS3wnSNk3gmDC27Y4YLQBYHvn9yDYs5o5gxm1MuhQ
cGHuy4lFRoAQuDtAW3bvuqgdFH1Tjq0OOo3myJ+wKnRrGdZpFBhhyy1l60Yob0O77izGay6FCOhA
3ZEWd5sYvWKiqE9V9nJ9c+UF1GnoxJun4W54nWLYjV9Z1ulA6LENWCfEJQh0v3llpLqNTdQ9e8k4
wMnUbXTVCoU6M0K/NBpipO5GYVXmapMAnzt0Mp0FwpBSLnfCJHktZLUTcNM7UsxzJgI6EL79W+OO
UmFk8+iQ0W3mj1JeOXU9x5iRjsTA6q4dZ202c6EiZjGFx0xA6L+2b3PsyqhfOtiIWEdwGDHI9GeT
bPujNp0fTKDJBOzuEPas3y0TSo1lBcb8siM0z52KInV+NVmRGutZt5cA/HsxeTfIh13gXF5itKwx
9t5ukYU33FKG5u4SDHDpc76AJ2CpcIS3lwbWtSrPTiSaMNf91aksBxVEpNppeL5sE7+mtgfCERWX
EeOTT8wANZGEN4MUl+nMtq3/HzWmKNUQqR9PsPy2wiQYihmppiVEz7pe4WvamzEc/LDaGTW/B/mU
IRgkRlLuTX1O9X4KPvbPU8yf2QIKihHAjkEK0/G4po7JGMBtVcI8vEzM4kacXRYqLDmTi9cKTTbV
7eHBLbQGE8O/k9WlCYByWboBh7CWnj1qMPuNjQzCfZFjTNR7ZZEcvaU4Dy7Tk+vZozantA2mYyGG
ggn+Qksm9po4K1aWzc+ZoHif8BEWpm/bgXBrHbw5X/hA7LqUY2x85OqYFt+ICrolZUqp4nqubsCm
FEw6gBzBkTyQfekO2FihIf2YP39jOObL3Q8NnVuCYhHXqYpWEdXFRFznp2FoSkTadTiMGB+Bea+7
zhJduotL8CaesdXCUBs3dhpMoQ46kAy1GnFnq4Gikuaa1ilFx+8nrBUxtyeY0jUrv6Vzosc3gQ+p
8pVTjBy/ACaW3oIKINapN7hLrQqwIv9uRQriztxmlgFlGXMrFoJxzimvMmCyQ0gGKpuJlWt7cfwS
gDLl0McW0KRehOH/OeK/XFFwSAXNTZfJ2xPJLKV4pw4zwuWsRcKziVeTYddUIYUg4/chOlaJGOZb
hyac9ysN5J8fue0wD9t9WLf6pAJ0a3JwZgA/sv5M55Vd/6RzzSXX8K1WwG4jYXa4SbAp+8r+u580
9dzJCZSYqxdwCoavxDbm4IPVkWjZHQcU2i7fVzqLmpkwSl7rTilberjSvNgQKpfHDD4UIrW25WDF
vk5nZg841fqPHmsLgC1wr6gAKrRHkZYV5A9ln+bVCJfgzjarXiasdFiRfqC4I7MQJxz79y7rrJIz
VOCvoUI738H4oNZAmNuJzruJabJrp5bwkGgKnS/HIX8gnShjMVrqRG8QeBv+lcK0PIuQk8d3FY8t
r9onWncMoAJazx3pmkkAsY+CBDCQtA0R2YZ0WpAVC8pUaLLmvzYWA90BgjvSiQngR/spew9TvKR9
SPIb9ZGybmYyByZQqYvnxMz8LhVI75Rx5VAtU+Hm1a7lxaJTmTrYfc/rH1e+9Xr0NBQhXS2uQzKF
rMVnMLmyiPZpz1owuN7ke8wNP5ijCdFO77essAZuaDGFXENe+J7HvtjC31u5H+68PASV9818SSIS
3qq0ivDEB8b18SxzqLPAKLIlNhVaTYWnSgr826Me0M5BOSyNU+QivzjUa3u6STXkx3eqYB+s+uPP
KoRVgauYA076rlf70WcHE8Dt+ARceRPwMfYNpuD/PLACAXOhyWr0cpjDEI+ZuJ1rHYTaYvw9dntj
zfMjDfWPrYWu7+J780i1S4ejguhL85FeZiEDrxzqyQussywHgAxr1CHt1dyYTE4Smwv+OvrD4pEa
wqXk6gPpKHrwTYGsARmmk3kxnvSLs/kK308ymF3ONqEHy/Pii/M6+DBglnKaOIpNtUwHUldmNK7V
CrqhykFqf4T1FKMTqriTlasY48c6IsP9oZcpbWQTQr0V1K4B4kAxgxkdWLq9Iw01OsPT0lCHfA8m
F6rwICcRbdTogfQo/acyWJUt1hPQqOHYc5wKdN4WtaMuroe7CEfxl1pAe8JPPNJ171OFSQ32akqi
QkQbJU2AhcueHxkpOWAhI65kP1M4yvb+mECBVANo+fhyPeeBAMz6L8N1+nAYfMA377a/ftN0Mv8c
srP8wiPExvUgTnoQRIm/szORP4pAUakCa3pr5TODISR1P0cLXAHJVN356ECdnD2ef4+GsrA1nABp
hyV6OZypWNt4sw/iU1OfN9A5pUbswbqHmvvkX3blIAtT58xHHIq2+5HZduwiwkOS6KnbNduF/fH1
0TA7KjjEoYl/PK1AsJWDg3oqa/A5a6deUdOwshTc6qA/0ctvLKMDaUBZtMTe4MXgkFGaeFCnqyKm
oWYmLy0+w4xiefclFoqeeQbTGoRUY+yxxhvJJToy4sPfnEGrDXVPZ/LM+kecSCYQ8+jSUohyiraE
ssZlfM5vFsXlhd1w3oCAF0tU6xMNcAzZZSLiKloJ/OfHeG3qTN58Yurukm1D+/PZFFHlnFQUkvJp
itv7zQd8ch0kxwwBPkigHuIrUhOeqbHelHRjtH51LpdASyThPqIB7wE0UZB9P3LxfUxalBKc8Q/E
L2c8gL4lK0gw9lr1oxBrVMg9/0r1x7E8f00WoiPxDvFwJNFBqHLDrf+ecbib0XVqkL9PdqUTrlwL
bJOrEp29FROyzb5YDtDS6qxhhNa55OgRt3qO28yD5SJ8Gr6tVQQ4KR/ZAaLBa52mO1qc2TcZjmgf
y348DFZcfZstxlkMQQGpg+kWHabDNwqB61CkoBntjQxZbHWErNluT/b49nhHDF+6wovKXm0GDLFH
jgQYT8PtY9L/DE++CvwJcr6FqL41ncZoQnmCTv1MDBNwPEb6029gOuCpPzx/qP95ZqUIoFeixYO5
RBeuUuunkwJBki7fD9s1E31pZDrcEp8t0zHb9jomflkUNj7rPVQiuy0YYQAwoiOoobfyacv1ZY/Z
66bZTrjkpein+1+QKyrrrzNH2rIHhpq316uop/+gQU9jID0QDVXeQd5H9UYcCDFdVNW+pKm3UxJ5
Z+eUrBn0dM3UXaPlP4XlUP8Sqh4kR/FVc1LmpN2dd7klmhn8ZPtSX53JXOiSz6smmh3MdWEW2+5l
97T2yoh09oTr47CafPJhVpZ7xHiJuplqYErBy+eCvVP8ZQ5OEZM3flfWE32kxzhQXwYZlz1eEipL
yAMALBTZSUt6wrFmB5duEmUF8YlvBfP0VLM/NKB43haQM7R2nhqD02XOhzE+VB11GR0scQuJ8e/x
ps8ZH3C4M6XmspNavWW1v9OcLjmQbx5q1mWWtTnZLz1CSR6CXYK5o6iNQEe+moQ5A8VKEHUaGwx8
6YzgnwK7bTn3vOtr0HhM7AIDEc4gmbxRDZ6OlDB80OsEP9EM8jSF3Nx2AOKtculJxno8CBe3LY30
m0fr3bjYg49m66RjoDAFcR53cNdDY11myvuPgmje7D1mTfIhAhnmURkL9bwHOiRKg4bvOKrQAcpM
3MuB0bU0wOP8rJUJKkQbJZfOMIEja/VNFyo6LSVh0SYvA5j0iUyGquQYvSauY2qFlxckOjpt//y5
GxRtf1czKoBTnG6H1IYLRHHudaxrPNx562EoyaGaC8tCzuW832jmHWjp3hQ0JBQBztFd37Gt1jMW
EGgKPCUOTyZ1aZh+E4lNiMmxlHHF6CdlBw5aINTvCfdiOhKIu2fuDUtCyaZrE2qtdV3qVT+aP2Pa
XTQcY3y4KSQvFCGNevxxFNiBAKFSBqCpPqfw88iHXCm+Jn/6ckaoNtcmkx1a9TQ0kDPJYV2yvUTF
6Z49QnGuUvR59S+Y878amI7L8A5EfBof9gC0WpkeKcJEldlL2suGb4X87l8wFUKAnCSxKvwlC+9D
F+6mbw6+IpsLzYgBRPld5b2Re4fkG0MPtr4do0rJMwtWoP9g2b0RdG1vTAlL2WFqB3rG+efyQIHf
dhpznscLPIWrEB/zDA5AM1IVEEQLrGGmWEtwiKmeCVHmoGlQJWoMzJ1YDydFnXZ5599t1OczZZVQ
bznG7pnHB8AwBN1rBnxm5BhvO9KxPmSdglQoUYlkp95C6TJSSo4HVBrn2cx5GhR2H9MMBuN/jqJX
U15hJLi3MH3kawNGppSBgs6z73B+EDynAxY26EWX0vEoqHmK69oEVFMKbgy1x2lO9YLv87vj2sFs
5SJFFzOaYhECBKMDqc7pKxmV4Tc52WfSZmg19d81t9edKDr52kbEq803aH0FWERoJTg6kD4IWgBO
lpn/iMMUizd01mFSUzhGBn/FKtdV/V5SrWAIYTmPzC/3TnmCELEO+xMS7JkrwR+iZb7/LxCqpEdD
6fWeq1oLpCOB8vbjfxGVC5BCGThjuLRx3SCTfbrroCUQYmN3cne/aVDtMMGIF3CVk9iZYV0ml5xP
HScyWIZZgJZk9Smac+RJaO4bnYn3LP135p0tYQxpMhjbHAHYQmgMk7+H2OgJUpN0p/hvIXvI9Y7H
Xk36+RKH6j6ALZSJYm/M0Atd6xOqb/wESbjjtDwHrxfRMPXUKJ7Yb7tPRlEunwUav4Ple/4Oqh1Z
YyyAx6ZdIn3YH4UWc+CcnWptsahLdsew3XVPGQ==
`protect end_protected
