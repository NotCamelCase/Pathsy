`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Ve+pTfJO0tadFKJ8MjNpIU7YVZu02So0jxTOKSV/YcPbZYf+TebheV1DKKgBOtV0vRqZH+gJT+DN
iZf1N+9hbg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
dldunNGnuyHIT0OzIGuU6yyNNWgituBYgFmMPzcj17UPyHVsgVw+NCP8cr7kiAua32A/xJM2fCy9
v/IjAnDhwqJ1kT/7SPryUAvmrjQflhjR/HjZn2CLeeMWnmlIv7c+UMm/c+8kqEur5yoQAOileFKn
OdLOP0cTAW3fi1VuCpQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
km9KWuaKxsm5K/650wA7g1a3nE+6O5pBCgfJCQRmvvkBXgKJWPC7x3MTqCM1naWUVR8C9OawZuNb
yracjGtjHiJPgSVfOa3/iBujlUoON3kMv1XW48KS4N7ti0sE47UfE3CGIYO7JuG9G7j17m4SijsZ
Ygu36g1JcseReeJ9HWdF/dvsGqIL/U6Y4+tJV+sf/nvWHNhjRhW9JsDQC/VLGJjagV90apuReUjF
oA+Wt8PDNDcWlCjhXO4wALLyQxje02buu7YnFDmThLODea1B6mZg+jqcHZYVuvgoWp9/3fnLOdjY
jdpwEStoGLMriZoNQ+615t3hztg6RVNp7iVpvA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KVmhBjX0TcPGu6UeXWAiYdedVkniLMA7e7JViG7vG+blt23yx2BwlGABWYs++YeMJNQ6bVfdZf7a
zdpIUkMagKukGmai35zLf2//3JN4MKQZrw3C8HUtmlK7BncqDMxqLj/ix0ExcE7RZDk2LJhn1wR9
EJjd36ksOVUWG8Neqg7S0jLYz0JGMGrX+mcWY2q9LLEpiFiSn6LMaBIjfwSHGHdY+Dj0ncVEtZLm
8xVD0zLx7JJujBUWf6wGKWv/FHS1iC4ZuGm9WLOuesBjeQit6W52VKCEkosdH5FnzpFOO0QkOw11
lkTYz+qPHi0IafEy0Jf+T3/5GIButax0qju0sg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
eYQbdhd3Le7t9oBpS/sq9pybMFcGoh7sezZQF6kMymCa3v99LgHRw9Al/WnegGrUPXc2NYbZIfqO
bbmYYHU/QMTFw0EjzrcwIjzAKPf7H3+OpyQ3nQEIjaYSSCZRIFwtwn7V2HeFtfY0haGSxHYZOKdR
KSxlRAehI0ZRWaDem7Q=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
muG28kv4DfheIQUHhdSWCZKS3Zl41dPzs/oR2ypUkxx1R7NBskV9CnkxPE0yZGpvMtBvtekQhq6T
eMZkDsigv/fEDGDHO5x4w1xCA6afVNeIJ8hqZOg3bSMtejPHWfujxDfEqU3r3eRWfctqM4+6Zzgv
OYCoqnVk3OadQcREDczV3FzVtfbe8GGQ5uim9n5wgVSzrDW/rRGOCrE6piSYN66qB6yutdYN2JlO
AHYNA1t8rLk3ykiriawAnHPnB+XzFuPI+Yc9wUYxzwKpzlW55d+R7ywDlcrHxt/PM3x/DTfZV4a9
/7BGDmYB9bXYVZ7BCn+wyU1YLkCGK7UpuBKQHg==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
lqGjHgFdU+h8voIhBAchHhvI4kbhE/DdAwRConrNorENDaDIdPwTK/GORNQ/p/wDtY2IuvqYiOSd
d+IL2xSkqtYXEaMGMkcPAnBu8BxbJKKyCplGiHrniTygZhzRAPQsV+MRWv/7B8w+bdfpKWVq0xWs
uBKjEOBal80B8jlzbtI48rYvf3o5eznAypE1UCtaaLx4TWmcXTwBgDfYRSuIvv/liMLpsZOsqPHg
T16FlVAkDSuOaoU0nCY0LD4lrnVFC3L7Qn5gHWNt7yIPiVxEnJ41DR4ouXIkHPz2LFkvRDQfJjik
GPum+ireuP8Hm9Pdp+CeNzYoXXmZh05SX8c7XQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DW91mt5eJqQ5mCzgO2eCAdTvNsr2FsfhZmASAubEXINV3Hhmx/m8ccKyScar9qy9gsbipQ3TKEO8
CcGqLHjGj7k8uFnFvM+0MGOfutlKkx9SJVIi6bK9sIjAPWDDOecyPEPSLaCf6SVoAVp7CyyMU/ZA
U99aHxRWqRUo2Vkw3O9hHZ8AVnxhiZivUpq9hYqxTKnBQuvwBfJIld2FYQMwXOD4EbwUzPDbUt16
O15e0pHxwVrbBSBjTLxWo8MUGWBRXSyOy+0Be061Lv2ShvsHgXUrhNeZiGC73HZBpdcTmWbOHVjC
8vXFgWGjw8R0rYLxTMJ6PNIaaCbrJeq+e8l/CQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nLze9FYLM5vy7BBk75IgxGQ43ipl/DQsh0PZz1L4XG4VgshhUHNr+WxIO47tLFDBBhTuhDcxvgpk
G9M+yzVDMmbrDvlEkj0WeN7V8VhHslT7FW8+D/mF23kgj5U9Eem8j17E9BBtV0H/PLJa4w9zsu7N
WHaNIPBe3sMyaYFBcLmRuFcHACnVGRJkLfta0ueiB8KaR9DMNwmumiiGPi35SUipcRyfdizO9+DX
BMouWewtB66DymEC2luKvtdnzVAqYqXyoLFkozepR8XgTDHMQURfFcZFfFCBpWLy95YJku19urRN
8XOXJhEnjHvdaVkNimANe4RM/oV24wlGSKx0tQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432800)
`protect data_block
E1GYftOMRZbm3faFN7gRTjrKbsM4TaYsBLsSI/X2cICy5PWScEM6+wvE7yu724HrpUnASNlQfitT
Yp4rThX6iO6HTiTYPsheqUrnWlZVPCD7eY9Iax1ZfGOcB6ZPA/UU1Gzf+2FB3ztCdERN92EPMRVI
sgmw/2kgsp8/JqodDa3nRj5wW1bTAh/+q4rHB+uPgohf8fpLph6uMkVILU+2GbSRLczhucyKw5Tm
U8av/tHhyTMd+5q4Pi/LE3tg16mHoSAF04E1bavszTtDnBK4pfwsoXvj1/cjU/KTeUoUfjYf6OyZ
tZZ9s4gozv8HlpTKmfU6lULoVKbghsq3BC3iXzUlDAR+TyFOiJlpFvg4TE9PCRCjI7ni5yzKXtAG
f7WL74VyJDk9scpZYa5QwJugO++za+ngFkmEnFuroPQLKcG7+1eHQjlOhF2y7R0nXG7ORitvnjmz
tVQFb0XyUAJ+rLD6OH2xyD/YH1tl/MrRAwclm+PkY9v3WoDgDM6acnbrn5+huIav3OoMa0utwYNi
9kqAD/5cMGb8j2NzfmJ3sTZd3nWoZjx/fMo1s8UPRT6lfx/lGRpw3lOvoRHRd0YEex2TiEbqFhuH
jSJfT8vjzdUhUn7ehuVhypidiC5s+Ud7ReGsRqmBty0ZB1PfR14gWSx2kR1GsJ2KrSQpbgZGOHpw
ZSuKIrwFNkb6eBz3mnSmKVxgkQqo1LOomjO0KHnypRZ2pSaBBBleXExtHWssyFd/uGERJX+XczXk
STeKIIsHeFnNFO/ceIJvUan/g1YxhdmgkXTvhwqlCScNMawGxebd1A3vOULJssIFfJ3+YQnvWkWa
TlJfEOjEBGlNECUXoFIUpzHvxFak9sQe3BnUvHriasG4G/M7CPpS/bq8ctp7w42A8WK4PCN/3Et8
m5wv74DxphNkn0//yyel6McigefbvU28K814wZ9XUIUMT5G/TuB9+XZk4QziJw77c2lVvM+eG2NC
gdlqYv+sfppot1kzbNhbrbX9YKs3cx2b4nlVwRvvzZKkCICQzmVtCKKDbGS/haDTwS9j753d9Cwr
FMeBLlwbuZJWyybRMru/4wmvJhfOQn6mh0F4CVgV5ZPoQAzvHvFcvGp7l9+ig3YHzMcxKDmbzcK4
lWwxH9xZRPCnOKMFDCecSHmnLcVkg9S8ROsLol1SzuIY1l1BHJVzoEj+OJAKWYodH5gSxugprF0k
qTMXly/BkdlmLj76LlxHMnPN5FtOw1/0j0pptxvPWu/akRw8s/aDtYhsjURVJEaMJyyYr1Y2X4ad
nNFNNeKMkq2N2h9Vlwtik4IlcuPmeEAcCdb1lFX9LqVGWoLktdQAuUWCVIFnI1c/mvieisvT8fTq
23w7nIjaTBPniTZ9JPuSNzIFLNSvuByK4sZXrI/zsNBncNRInEbptnLoprJmtxKe/5XRIKfNbmDv
PTo9UCPWZYoQpzuiPfQZmjRVQbQnu0P96s2PneJ0ndVc3rumz8bE3kpfvU/LuIpoFwk3wJ7YCKfy
0QMDsG1cvj4pHhUL2FSzKx4YiOwGX3Lt5frHcC9kNgxWJJYZxX1GWWmvAwlJFnpUBOwrXzV253F/
meUm+ubYo5uWIL+ZLU2ki2WrRqhjLTjQxWuBLOywP36YoSvXFdsUspPKifnvQsXEY53lXTcFlMOP
GR53KK1e8eaH9tSGrZ7uwWy0mNaLy/dh1Ik7Wr8oSH09gX++LORPVI8CDu6qT+b6iw0V274Zmx7q
SM2xyZXKKn/62MX9cuvzbYh+dwXxiXJCyyEzopDT1OzBtOuZrpy0tniYko3GZfNv494aASrI+3OV
gGCFIHW2qigBVTW3QKlEt1/AW8dbCosDbAWPC0HnG90fTcrjzxXekytXJxbDnGc5j7mRCV+YgBDD
yRmyPJrnnG58FOpeoiooNY+e3zlI06/L/uayn4GM+RZ9aBDdtiLJLpmnxkrDrfoedP/Vk6Znfv30
xVfyVA49IMJgNFHMJ4JfnM9oa74WozKqd9mwMOLDNG/84CpcoByal2nqn1yXEMGAD/W54Rudmf3B
sOlXAANvgHFmc/xmia77aoaTuxF3HOZl1xHXSteB9z+Y3tYsgbqK6Xkxs1wHnnXhL+F5LgSUvLQK
JwX0872oQY5Kgpk/yAvHXYoRujFQ5RBKmn8VUT/EKY2e9fMSfk1x/PdxQ/nIg/p42Wfy61ImV49M
UjQ1g4THJ+KMVZdCEIP88hM/eKx4cSqT55XdCCGpfZ7UBcHmC93UFRRL8NVAoebzG6oqTqxaqW5z
hYslK8xjrr77c4XvRo1QyearRMH04pX7wjoty0XkG44wxzJNIqV0/7liBfj3quuMo9tSBUh6OJG8
4T361DLFDQbBQeJqLSny5E8OZ1rIUkyi3OFdNiD5gpjoWPcTVfW4hCNXbw2i4Hr8qKengbpyYI10
frHMuyEVwnmXGIaodoyHHS43osJBP/T4IjoioezwQStr1gBnYwtAVVTHaq6ZQWC9ZNNFomi70iND
idiug0tCZZOGkTMy3ASdPFrwWe4Ls2TfHtq3XH30X8a7WC6eK9JV0TkprIbRbe2McLl5KwM4eS6r
XXsYTd2SA3NqS3i3uU03Z74JS+gRgniYduXfVHro028Dm1peyxwtk6uMfP2KumsdRtGkYxAO3x0g
BqMO8H1X/mSJO74zjR5+2nYh1ylyO6Y2s/C26FebTbprnUQ6SsPrmigU0rxkcLpDOE9iKC/zPxti
FyRRbVWuMD9h+2PRmOyvoU9XXMpL5uVq5UQl5EdWgo9nt348AtisVb8dwzCBcC7DM2JxABVUtK4+
uqq6Vo21TdDkEdPjHW0aeyqvSfvyefOPxz7sEyDeK4fZeSSPIqdI9OF6yEt+jBZglHB2TC7rOEKk
Ht8VQbmkQrrqxiBlscP0ndkkC5g3LN9ADpZyThycj0Bgpo0zrQiV3E3ejEL/TTJP19zq2gQsdKh1
78B7HRyijMOg5qLxPF9c78DdPfO8xHV+lni15VQqv55mBVM3veFQsKFxDPAo1orDOauWW686zLjV
SKZ9ncADkZqTn8mp7Kxtw7HMZixi4NMGx4m7uDNH4R7VtCY1DEvfFWXgnoRzPeEGeQVFsf/kbND/
POHGWOQGxoqHxYBVbbxZQfXMt3EsvTuX/OUq9tqYVm0Aw83bhp6vprdXurpXv28pCwSMYUAvVnkv
JE8NAkdTmkjOWQhV/nDg1tpeU7gp+vLOK/GbZ/eUUCYH6nWBbOgQIJkiF1AYAZ1HSot8G5bsSJpV
gvFqtQv8p7yiphf7t3MzK1sWo0rzIYSjvqFEeEQDZxW2KzKHANTlF1vafEyUQjgKdBgf7XBiBYAp
bVTuUtPC4XiQQDmYOcc3CiJ55+PKOJEtyQ+d/R2qN4gNwB3ghHu290GdXItwrNDAfPgcdqTXrDFm
mxd1ZI8Hgzg2w9a3ebqMiMvOdu/lF04xwyqyDbVd4n6rEql6A9fa5uU090WYW1ZU2++9YNZ53N/Q
LNJWOELIK4Xpp9HMTQ9S3/oE8ODePT025KzAgC8mCfl7R2ZyhXv+yB8pCycxz/mYTNvaMFqEP/G6
N0JjSHinh3u046+r+k3emWGYHItcvqAuZZNQEAvijGiVi3cU34MspcYGfnysXHo4Gw61swTdQMnC
zL9rYkCBmosCLyly07u3d0+xoB9xa2ohZsP3R7kKFrwsc43R9dURLosLOmhLt9X5ngfqWi60GEAx
9iguqLH7cn7oSKbfWwWIodXChXSrJ8Ykp5FIJELIYPgDpGCJ68EPpDkAJV2xy5GBWPkb2nj6MC22
DtmESPeUsp2m7w9sRAkr6jQjRLZBwTRJmByDkpKx2ACfnsBiE1M+K2ojEf9e7UEQIlr1PcAZ4x8w
KOrQx4Kx77jylaZyh8MgFRrm0+QGalMxM0YcJ0b5Uvl+ZwufEIhzerLKnEyb6QxI2J9i9VV9ZlPk
WvnGqMe1f5fb3KF/Y1omxO48wYBd+ZFvLgWIgMhtLWojHq+qvf8ExoALTeMgSeueGSU5iPqATHJT
ozFr1KvMWQMz7fUVVmgDa8lOJ/zVdv4vTTCZVEsX1nPRZ6b9PQyb68nA/T9T2AmwlbInV+lmjd5b
JR/plI98EbMvutGpNRpNFyXsZU0R2vaDaii2cZujYFv7GNmCGbYvgomOF/pGGB7aNWftxsj99ip3
onwswqCYHXbtWbHxkDI+9dvVoRUmHT1FXhT0facbUJcGR5018Xx0bd37szL1F17ThGD4qyeE4vvX
olkt6MOPecPT8XmojrZrsP/KLut9s8jWMArmjic+cwVN1oaGdakRXFbGDgJ4ZOpvq2RQg1DCJ6y9
/YBCHLyHeq2I24JSZBaV/xSBu2fwYy8IjStaOvmrKChT+yV3XQ5/TFfBQ2G8syEKzMz+gi5kBKck
eVgPGwOlc98oEkfEP+60GR1cqD+xSLW0jadCXfCO1jN0xEhqr1exW8zc5DKszD7ZEMRWB58wGl/r
ETFDGC7/ZWbLGTYZwmea//MdU+tkmIp3qUnSS2luHG4ppDsmX1SfVnDFNuqdyTLv2HCI8Mpi2xqc
AYEET64DzeCHjluMvIbqo8HSQHN5N4fkrZT+u0ZFYZv2tAnMfpeVm+DnCECYFCD11C3794u0B16x
hNW/I8CYvrYZv1D3rIeI3KEvRLkUKj0FS16Xx48YoDQ7eObk1oiyxa7t9GuLH62ZQTXFvf0kUJBs
HuAZfRCXRKpwkbOR1y+XKdsSEJwmH9eB7SHC4Ly3BiUNIeQiaRUTPEZ48gisndS4ruQrRoUR0xep
Blw+Qg2jHI9Ri5b1XdtO46wdoIankq1MUaKA5zmK63c91Wv9A/XM5mnLaryeiOM+sg0seFJhUxdK
GIPmtDzi+ZNMmriiwC94OECDkikHzlww2p501d8IwvFlD1JPUDk8VyASPNc4UB8HypSh7wRXl3Ol
C6kNpZ/oxTgPSQtTvrStnOK6q6Gq53ZjejcWi1y41wguZ1hmgxFoOw7hYYRSM3qlQxogSy2Ffgj2
wOxTFmle2mgaLr+CO0wk/0rZ8305OL9G9CNclJMO6blAvviviLfXZg++WFvHw23gCwTyZ9wKiDAE
0ecNeBskU+NT0A96POo8ehHy90q7o/rwUYCiuBhJXFkV5RMQqIrU2DRkho88y1uoc4C8Nu28IeTW
z6j0m+PKP5bsQ5uL7+lLxp/4NM//kh1YJH1QB2olh/C9/p3GpkNSykkiI05LEU1xRCBZnGpeOt2x
PFLE2wEK3JQteXEYgBrZ8IxJ2jJvFqEUeWTUg/N34lNDcTGdpF9rw42Zq3mi6lfefiDnfsVRqXO9
0cXAA3e5/sMz+NhdOq1B4H8z22qvRQsmg9mymSLi+41hp+yo3r2Gob3WLLCQGTpJ3zupw0M4cY9Z
DEMCgzwSMAFXwomNWHstUbehGUzgiTnYlFYGcpNYMhpG1RsXhmBzgmMcHEvq+j/2ltPr08mWHLnF
TM6lnpB2oEgpvTTzlzc6XskBNIKPTY669/c5wxvjfKrcowehh3/X2ZISbIMfiGHx/BJcvw6jZ28r
CvitL9qs9aNU8s9CmaIv2oqRJBnOkspfewVuzic6v6Gz2HR0RKuV4qNeDKSFKYy59PTfEbr1MMfx
YDTGP//JD65TD5HsdOT5fuz+YG5+R3gw0SPEtKc5UcFI8xz6NImrRfjER8vda5kLMvjJ+zKsnwui
nWYKFjhpPzciHkAv9KzTdS2yWLLbGgMrjxRcjw53dS2Fz3H8ucgj97hRAiTPwhpVZrg+20b2V5Kc
J+LLqs90P6VBWbY0uKKm2WxGFtyFYc9AqNTdfwGNYScv/sHfp6zDKuIVpiXEaSiqxFsZzA+gKaB8
PgRfWYUgcCVIEQXkC0Z2Xn84zqbyzpwiRGqOUX28qqG/wfLOuB1+OZWw82YR+F7OiZyC7wgWuDk1
QoGL8iV4effGcD5/R7VR4oBNCZLXo6n1kqpqqGlrBkl6Fw+uWnkR0BwlmmjR9GiPDE/Z3inMHwl3
8v1oaRlmm+93/zPqvdCd2wzacuXxkLaL4rKzemAYz/8qCLCFZ608RQcCDTdkjyI4SEl63pRYJTZ0
amEJeFjsF0FCRvledO/uxN4eXDVtN2vRIxCgenfqw1VwM4yAUXKtA4DiLbis9pn1f0Jw+XH65fv9
MONc5GbRb8ItjJ4xiU+KC0nZ8kfylJ1eDk3+096JZSjrlz8KS2jVV7aM8KeYsoOUREK949dsIdFm
SAD6YfUsRM2CL1EukTWSsI+YMeVmXi0deMoQpKC6rgbwEQAUL1MrK0SF7ceC3jLlHEpGyLcTtHJH
qslFvd9ED+Aly2P5OLQOkD3JFl+hTLEDrriGasK3clYPZmvP9aIaUqoOuMLloyPeBtAWijqUXnG7
4GpWIhng/KVhLRKCpNvDX4Tw695VUnIo0wx1OH2ylZeX/ENIGoaRCZkpVZLReakMR5bqnfsoEafl
vxHnacPGVfu+yBv4DUOWxi4mxkvRMYXA19ul1egwywFj18XWadhari7V7SFUbO3aCfo04auK/acS
zBdjrmBwP0b3lCQyD4Dgq/iEnIhDdFopSJW3L35y+8FUyME7qDjD6zVk8Mo1OP4FJNYD5b4lnibH
z5gX21cVrUvuscXiUBAOJ3TzSdLqUzwQ9b+ogZ+hPH8J8wXTbQqVikbx/eFB53SZnj5ojmKFBqXb
dX7lkM9eu6pYmrY89A9tHoIL8Bp32mkqGHUHxq/dIiiRI7zN3gMBoZNgDTFnfnockceN8vRFYqCb
hT0fjU6Zt3JAwHIbt2OPj4/S1PfEQ4kegddAeIk6aqiCfiIYoY25CuAwZzsJblECiZZ9ua9jK0a2
yoqNfHXdDfqTW8CW+aI3jhq2I6FInomicO87hgid1buNLntRpMgKRN3w0V38cxAVg1pptb1I8sHc
E5EyxzqjnLZhWw1iCVDUGm8kxlrKeG6kuqIA/eVHHIvNY3UuIPkEA1cGmIWyMytdT2nK8wcUKDfj
h1pOKNCF/rluGj4reCyrx4eIpF4wbH8S5jYntHQpsY412otU1jGriVICw6uI7iXWMFcrGtcKL17A
uBU3yyBQOxtohtxEihUcTXPBaOTIJCwvGwxbquyYeRIcZMSQyoDSJo+l10kngmxjgA9PhcQ24gbJ
lllkJivHdjvEUp8XDmFgeskyJtMDlWHKWXdwXibkN68r3vKM6OQLSJa1n5pB1CFjwQYf1levexs+
QxCTA3G50QZWDFoStJdJUslhf68LpYhp6lZiyfNCVOoe9m2jwO9+MfISU6dShcwJM7r7Jg3kZyI7
uwr1up99wpu8khzr+8tSHO3yoSJclkU502Ix72BIIwUkbvHT/em+w2kx4btcQrb3gd8wDZLOUDtv
8fXHkd2W4IH8on3Esi0LMLp4LhK06vTy/UKaeY9ZF6QUC+ju3pkVB0wJTsp7Ks7sIVGHleRB7i0d
fzyO3fRR9NTOSh3txc20B3duNQ7ML+S8BlryYBOlAA+Ltawe3cUdj6MYH6x4fchX96V9I/rQFyrt
5GWMlYPnrYieNjiLEZxq4CQQu50odyKHwxrb7GDuUkvHeqV1D/tKKtyZeyYeQINSQ/pqFV8IwRZF
zros8cP6g1fKzAwHjoKWi77Z82vCDZt3zUz2jZ0PNFbYcbizauO14cSt9Ec5B7XkMCHCGPWYdgnj
lHqJ7yoHbXNyU44ljIjmihvqfHDeUbmySoFuXZgOnR2CQ+XxvdjhTIyt+qYzZdI4hZFEZKd+JvHj
YseIUAKbkgqg6iMLiY7KFwgXxKXege8SZFhACUupaxBVYu+zq173oOMbYFkJjv9MLkJg+qrlsEn6
hBjz4kNmgTqzjLS6Me2AgZNiWitonTj8kqUe44tAFcFHPFJycpYuU4ZF3buduz5gYOfl3FDPjsmc
ycuLoJ30thYnzZBRaRPec0m6r5xe+px7POhGAc3dLTWTNjorvzScNBMywHe0A4q8cJwB6UCkS4C0
3foic7TnG+AKwrGw+XGrJ86cbi1YFGko3sh8opLk3o3TY7AbqnTSM5N9jwQOHKsB9PxH0+hhBD10
kYF5CFxnfcS4sSvs238SRWgJmWne2W1wD3r2aezdVH8vCx2JW8dxO4Wixa3ePUFnFqcXZ4D3ov4v
7mBgSlTkFbkl1Tt76qCn6X00HM1RHKBsWhzvSKAY6b6rJLSmz8nAjiD67IZDot2mAh3xJiBQDUkt
aMbFQRbSrN+vB2CgIxsN/Sa0myfCzSpvUt0K6X412KLpTCK8ihBMxdP4lC1k1M8DdoV5T0676PJV
AAA6UemwyV9P5IDh+wZAV9TCRtShW/QGUPCm4bbuEcY6o8vGQkQNv6jq9ciR7UqDiJ9Fja/nnCYB
YgXsAd8AY+hEtX1c4Le98+Gein2feKRunN9OYtWzaRNju7oHRhke5w/hQ4T+UnMX3u1JlSLEkx/4
8WD33c3BNAL++563AuaBM0t3v440vyeZpK6etHs18+DL9jEBfISWYMx6dBbiTwTlffkf+3X4Y/uM
zOhqYL6rxqzxrd/xudfKwJmJpvqwNWWcEyN2jurtyQWOx8+wW2zgskNn7wa8hTg44K9TTLyDU4tO
4fewPSMvjuTW+eY6AICc7ek6lGeZFvZBbdAelrXOXvtp7D36fn5BOO+q6IZUUdS/dn44plo+14yq
hFRKsdvFnBHcUW9pceLx1Eb5mXSur+k94YMTJlLTLinyEJ61ijYqbOYzElPQueiUpUZ/eeUI2oYy
QjoaAR0CUPPjk3Ag/hCWhDftyof01qCUTSUk6PBlQBcayfsoep8LXqwCasNuppkJXuitn2g+Fop6
bh/3RG+pe0rL+4lgzDhjrtnn7TO0oGTHQMeP/wqsLIcMxfYpJk0nM1lSCsml8JahD+wJtDVTrf5V
vExkg13SnQGOezlP4mQ7MGMcqrYepCoThE7bCzRekYGFMCYUhwYF81hNv1gGga27h2pgxBIcHOGj
bRJW2jRB/Re7rEqs+su4hDWwye8n7SZ+3L/2FGUGOSa2s8Pk1ZpefLy5I6o3U8PBCpY+Hs/jwjlP
20BpVghrmwDxs0NtNEz88t2O1MtgiQwcJKzyGZp+fJwU2DQ+XYMHZLTxBkFhuX3I6ZzAg8ldy0/L
q+wvM6ZHUKURSDfhmD0Jjb1s7I5ix6+39XaLVjA99KQqYfIEdXuEGl2SGIlmEEic1IxH01k3Pg1m
35eJdoCEbRfvOWAyzB08olwn53ZzDVpSfa8sW7a3LhjIecKwJwBFsBh2mDhhZMr6ntdT33eGl6BV
u1VJ8FbLVfccud+TeNN470R8IvC6m1w5CFCAW3Rl2TT+kWAEABxX4jdc9hhnJCkaf1geRYPbw7IL
WjDSCZZ7qiiZYZtfZtIIO9P8qkGDUCsdiSK/8GFbDrQ3tx0yD4gcE6Z15PLcUVSLVqT3B4mL4k5X
xD3GTn/9Ybbuksh4X0wk6fIKv14p8ZtFj/6JDxkbOBsbn6mWbksmdIZRVxQ5ySu5WrhbCFpbl0qr
hahRwjiHNJ7ajwBysAMkF3EqhdxExQS0nRjrG5MutgHQenUfNEUKIDmBeNo59CirDXjsDDbRsd4x
ZWKwqk0xz83Vo1anCbXWqzTvna3ut/tAmtokwcCuws0MRujYVuqlGQQTtCm67fUdf8ccm+mcF4Cp
MPzg8Y2sDuvCa5YDaFjKEyXrfS3+ugZNHD85jh+swrCRbxYOhO+0e61Rz2WFJeBRbBI7JQ+hj4td
sL2mTiiIZU7vRMI1xNEpMUkuyw14PLN0gytFXK1VnTgMSkxMAKk6IIaMMVn68aNVKBpu98OYm7XI
dDqaD+5yeQBL1OgSQ2i+edbRNGsijpwOohXeV5dHgxJ7EWfVsBqNHcf1TDsurwofqH+fkIUeY3tN
M1o88jc/wtrJlodZYOk1CP4GyHTASkhXj/tvchSBlQjxfQBAc+PiUpEpTNW2MgBS9U87QR6SxATc
yBkTu3viHGbfOkjjLIbErYY1eba7AEIkzaRjjMFR80G9HSp/4izK7GOXkl8IQc4HbeAkj4OU+uJO
xVut6bcJ6EYGaexBJ6NJ+MaLfEi6V0f0+/OO5too2fGN2ByXYDOKXB6g+KJp1ir9NFMb8KlRpy+n
MB/J57KbWExOuiK+NAX0TkBx6EWFbVoTaalAsDXyGm98baFbfJdSAsNsDCPlVV+ybYsrQBCVUz6q
rjT9bEKTVxp8kk7giouxwmPRLzuGPpMOE07+uqyE3ASRrRmPTLhGNvyTqpGw5r8kvv/n/jo7kWZY
XEO0WpEuJZC/3Ezrd3NlOGQs0v4tmj6BW+hoabd9LYNVPnlal7YPKPa+76K5lFJkPpSbSJGCeDVh
RC4ewWC+UtyCbLIZoj57PTleUn6qPkhs3yLMOyp1xVW1BVy6mgluVM4bDzPGveRc5tncSgFMXiJ4
tQiK0jwJP90TARTHLPzIjTkUr9GENOhOUp5+Wz9N8+mUyb37PYPFx41YWQeltWCNjJWBjbEEx85o
X6NRrWX1DGOi+iR6sWc83eHVCIxc27POSPdu28KOUkW15tmhSVr8/WaXzVvLYt37DGBRqPTyMW+y
jL/da4iYdiay6MZH92SIhEKpHBSwBR19r7EDLP5/oHSOsCWQS5z6/arwq2wTcwAU//A/zoz7mOEG
JJ6vYIXE9VHjbIEwxS38K+H4xs/kw7vu3baTNzL27yiACffJTLXlHUgB2Ly7+yES2dAfwlVX4nnI
dAY9u7FiHjRojpT7IV7Bw9QWkhV0881JZIQ34U9WwDuDJMD2L3mW9ZPoBugFuoXDSnIGx5/nTjFR
OIDPlDp+Nj5a/W+fg18QD5CYS3PC4AvO+lI//9WrEz+vc5b2HZQruwNR8yqgTPqyLqJ36ZH4lfko
BQGeePTK0qvIlFYTXqGKGIGDU8ULErYSszET/0pRxgolCZJN1hdl1sXhcNu6xvfUb/ZSHMCSYyyI
XLmjokS+KoNd8Hm+GV1rO4i8ZFfZqGzTCJIBz8qDxVUjibVLEVkimUogVwlOL4ZwVe3UAre37w5w
+cMZ+pzabCVFHF/RIAUS0M/EBwHGQEzO5TpjbEeitXJkmVE84aRTstYrHZLxH4ZGMwW2IM18F5/B
00vEB5Jld2pSc7U+dPgFM3isriko8ve+wUNp3K6EFtHbxuFWFAmeBxOl96oBuS7KRfmaoWZY8LSJ
cg0SkwVWYSJ021DLYa2Oj52wjswdC21jcRj6xAEpkCDqKCCsGirzADRW2Ht26QcfftB8zoj6Q+rh
wQSrExKPxlcoh7hcFK13yRFj3oQVhNf11izdgyL+okyFzcP+hhK2Ou8/EOhU2svE9lDF/vPvb0Yr
JKqHHqWM7uM2YoTNonhmmtBaE4T/QW2vyDSEgZGsfUouY0k7MPjR8AnQlnJHXBO05/J8fYxuHVy3
o2GJAyPYcD9lKuT8D8+346ohwxdgU/GZ8Sf1MpKEgtvGCOmi4tWPB0gP78jrBTctpVX1X0eIGAeh
HF0DPsc+NUXUAIfvc+sK7+A/8JurwLHuHO1e6TzQsc6a05isdpJspp4fxfuJvU0n8AeRhg7t6wSE
1jzJihLnlMfUpxsvr4vq1OSfvwTxqQi7i0ViO1B1h38llkXAqOKR/dHTSMbU2MC0XzWbk1vwgQ1G
xAcihkrXHcaMxcwNQMBB5YwyzawbiK0TyUz7KL6CzavbXjUm0eKyeST1S87D0hMkF+czBqGV91od
ZbzVTTlZIebKyHTOj2X7gFKdMDd0Xs0FAJuQvQlSybaphPQ/As0W7bNMtLPxZRR/E6pSJf06sZTo
q902vrnaBsLrmFlFu0XT01Yi+noNpJmazElK4yTS/DF1BqLIp4mg/zvRJAelS4K3GXhBmgZISIs/
e4zQDd7yYhxk08CClJVqhTaMj1Y6UpkTIQtDPSENrpDUwSq78OiNwADNI92m805VbkRs/2EsdBhn
eB5d7k2bSygED+cc3Sgsn6nGpdk/0PqH2hjNcWAW+w3yPZyvTd6sWpYrE5o7bXMbg3reLm08fpkc
IN7JTFS71p6HjPaxR6e2FVg2sYvxZSn4R2/BDeDHZhLHj4CKFVUwZStAb56+NIyh90XgUNODpTue
Res+cS8cP5h9GFqBQitVmBIPNr2ZMDs5Ak5X7zjsyIHMTVudirR+Qd2KoxAG2DbmG4VOqSXqwS6N
cRNkmh0n8qedD5RhrIwRvs0PD4mAWVGt0oVvFLs3ZipUeJkvB/RVxw/z+njoE6LN3eTpynZUpRFz
+snTaydZrueyzux8zjFsQfksczgIxtJeKslVtGo1wgq1UXser1YYrpRMKkc2WxtM86eGBF3Mjz9/
Knskjhr/J+jPK8nahdfpQB2fKVH2AZ5cgH+4uM85e/W6xY4zP+iNLVyYzzunFKbcVAEcgoQFT/7c
P3qILqOVSVnrZ8gDYxfrHEOzMn0gSGCdlTilA4ZJqE7SGs6TlccQYvfTizapzm4tgtioxKZQim1d
7Wv85EtZnKExCpKXcnhCEOH7YYAU84Bq7xcJih1W8yEbdBaRRspAyS1j5+VGc5J1Hyoac19QxEt3
Ft0dulGzalzX0hCL8RypePOQdbKRSI6YxVU9gIlGn2djexfYzFAHzDZt5acS6FrBZCqrBGbRpjNd
lv4Ft7oRzD4vQ0UmuzksSZ9fEzLFdVmu50j/gvPUN5vRiUyOKnSWliz3DQWOHiStAJqVmfVg+YM9
oFtNjIUw5UP/5cIL0LH1JsUkUHqwlyYi9TfWMi5WLYt1QO7Vt3FUrKSOK2oWO6g1nvLJhNffSVrX
ajO+6Gqza4/iog33L9mFArtkp1J7jUum8sYy3nGRD6+wPBZlYhSHd1J0qWBuFGwwbiJwQ5ZrbrhY
HEzeH3U91qvneeLV9S0iy9O/Gx24Lk0wBv6HObeGT8Qjrsu+11ofzQV9wjWtF80116yRwdCuXo6X
VGJKlDgCCN+WXV6Am6H5rMkAmbI+i3CpPwbir5q65FRqQYKeBNuZ+gNe2xQyr7P6I47mJhaGt2OQ
2lqIBRl1tzJeNBKjHj5dCcnG8iM+XmKjcJzloQr9IMe+OIZS/RIyJ1gziIlbuhNOkPKcHUQs/HuO
YgY5YexCi8yEa8P6dYlRBOuTso8JCRb2D6QUKuB4Zq7P3MF8nnJPMDV3GcJpKzybfefxglXIiQOp
00gdfkm3RB+vVyI5VYR5RHZYX9bnygPKNjvsZ/l4L1DM5mGcICuI+vRaBVeiqEiwqtYFrDi2bb1F
sMu/hE0mvd+aHbyBbEvHyh/vvgEVV10G4Z8yYOda99bn8u/rlj5axYkE1ciqV2bTeocDDreVyMqA
y00TK2enIj4XfBHQN4uXAL6BmYCLqqCz+DQpxfDh9dsTL3hHkrragTQBNnWEcE1kBAVIRZSsb/9l
EyC/xAeViV7uFwnbneZMSpQGzTlfycnXkNBOGeT++jbni6PC9C8GcIGN/t3lPlbKPacQXqKJgVwU
XolYAKHUN0rDKTWZLTtb1A46hKPnuBVNuIpR5rcXE+Hr9Y1K+kaKokDK/lStRS4dsT74d9Wy8k0B
5iFvhRyIGqmwWxzdv/nrSwGI23yXKiec8cMg6+/0cdwfnhugvBGygStJkOtk+PY3yCJCNLYfOtGz
aFbRgbFvFs03a69N0fdiQ7G0VkD61+0DiOzMU1mWQIYiVS9cvdUq/Z+SUnZ8CQO6neoDUIJI7VMA
S4wonbm0y3Hf/7XOVxlqs8CbR/78yILzSPFMnakuCJ0l4eiApDi/TvaMr4ayFqkGDxsKxAsvu8TK
kjTg4ma1/0Tkr1dJZbPeaWbJtejJ3ePe97jb6W7KHo4is1QYbAAqs5I7uA+nZLOE3zzmVi5J3euD
SY9rRcS1cTbN/iSXoiWvIPT+jwIk6aeDuvNfv2Z8M3zxipGzHJsQWlWu8RXbKT/zG8CSs6vRPEVw
0RBf/5EVj5K1ZbTpj+uXEDCRQJTsx6SW40gft5xGv1kCnrrIBke3OsDtGDJdX6RghS2iNSnEqf8v
+y9K38q4X8sYurpqndAr0HTT5HVTaBR9cKiUSjK356GkXJWrB6j/zreNrOZYzGD0A3P6+W2BBW6r
o6HbiyvHvqdYvNv1P37J7+bRU4yIm8vpsrUAsHhyyzbc6cxN1h2M1vjWhi0My2Ak5SxwLMOlG58l
4adYfUQfAQZGI2J3C4itN7+FnJ8wRfqhrmzhTvPAK4XquUKFzWx7yKBy9qf0N6gRp3/9jPSmYZaM
4b58ZKL2/aNSaK4Qf5xD+ETnZjnQNu0Q4qX6vcDhhVqUylBYYj5uB5gaTTD/UF3q+7m7yOJShX3/
R812XcyEcV//kWy/g8ZroujJR2gMH16he3znd0yIvHu4fiptCXxUly4A2vfiwFXMMDQJE+EidKOv
lkyLxuoU9fTgNJlE7o3i+arrcdKanQ+Fh76sQz6UDDOtUiLdkJMlO0vDVsI08/IuGMHjfwPzCIcH
qiyhylG0+MHh++BdQRyZYVDK4RRzpM+HvVVW3fkdvn9PUBJCGd87B+DSx6+G6lwL6l0KVtccP1wP
cOjOEy17guGvTfkxnocarGs7AqNPuzxKlnnmdqB5TEeIiTpaAqUE9BA2yNEH+xW5Xyp/jguSInQG
Q5sIrswMLE5tyBy5IpsaQwoNaGCL00TxDSohb5DoYOLwMEDku+ARiA6wix0xgoplEosFZsE4nQBs
4K6BTJqAb2voWOx9P9kGE0acjGqZZkEOIKC4qUnklsjuQjpaCtKyYqGooZH39qCrq/rrWYW4yJjs
//qaMnxLn4SswQQVYgdX406tYrf4CwPse8PFXb33LHfn/t8E6S5fjqiC2+qx5KUvTgQFTwPrsEqJ
/kJAS6p9qyI5PR5DWKpvQpzYC6qZEhrPWUT6Kh395gY7EMAedXkROXl4nJAF+bpy90C3AzuwDgEb
olXaLvNcUWeU+TQppFbQxjWIiOp+jVU2eJroq/ukU2Y0kYRAxNCBFcygy7+ZJdKkXUm7jSjFsDeo
ReDgaxqgAZgIz6wmFUYjmKbOxclPIYAor3foogURUZQHhuAg2ASZte0tiF61VmP/Ex1/bze47eCk
cijPVCfNHwdfqAJwMI+EvJtNOlkb+1RuhD+VWly7jNA6hUyjqjUCUu2g4ow9gEA2b85tvKzaIyu4
/pEpjUfVccjPDP6WVxZjYMmfGpMv9KUURFcjfnq2tNVj7anl4mJbSxXTUI+XIfU51czBaliqKnSe
g4qQzvBZdBhGjMcixKiht19PKUP40zowUkY3s/W8FnkcpChTPoMv9Uiuzi+dm3n8IyvJKuaRpwQQ
J1mxgxmW/JYfiskXrwuLi8lAbnRF0uEfJWG+MJLIV3P8RPB9WSkEzX1l8OhU3fcJpjynYouAD2N2
+zFcCVFsjNtpMn7VCB4l0uojw5WLd2qeUHKQJ1c6eUymrOPGhWGdR/FSmDHCSvQo5ABSr9Dztbkt
nTcF85H6EQ8+QHapH6v6iAwXRB+LaX1pKWw8metgAmDZ21BNr3ftNZsd8cG8nsnc3fVpKojZhEsr
JNLdwu8HRiPu3solHiQ5YJt0XCXP96MXv/8Wq1sDfxzTzDSHmHUIWQm4WsER0+9Z9uOQYBTUF64v
S/ZYPyOssukqxQ2ytFfe4fKDkzKp39o8rSx/wKwiZfaPeuUEMPRHmfcq4hfS7kugNl+rcv82H4qO
QfRGmMe0m2jXNcnzTTs/3xDKGQeGM5MV20oSHdj13vt+SxLAHd9TzKCPLc63YTH2bMTK4Ir7m/9N
2eEhfn7f313PJOISXdqpsRNgCE2IiMREWxWGu01C52B2jjVlqU0+qCg5gEGcqBKq1QwIqaZftgzM
8yDyOEP68ukPZRJ0yOknQsKtakSWmWR0QbKcFcGkJ/rVEl31Iwe/MspjtormjHHtLjK3BN1NjzDz
e38d+bRmzmyLLMAodyHE3DrFujC2MeUHYnc4FW6VRf+svaEKH2FFgpnqgMCASkPe1Qz6F2/eQrai
EyNAjpobHD6mqHCD/uv5Ni4jVvNGxSal9AGOhj1es9FV2qO8mWw8S6aIAxPVKzcNyzHYni+L49l9
cK+UIwAxAdr4Me2g0ThIqpZQeKXa9Dzn0SKeVBAUPcLykx1JzRPe2Op7YW8mhF6QoqwPQ3MRX4/1
OMiIO7HI0fU6mzFuiCNnouUv0b7O0xQ8BYShX6y3um6ot8q9cRlnftCBmYVAbODMBEfX8j8bUJQy
9QSgn/eoH/R7KjsFwf5kfFWIQniuwAVQaZPp0bnVm8SYmjYm7vOEjanb+es0WSURqGuI7OXPIRiD
UyjtyYpNBaJlrk36t2RhlfmrXerACrxkJJ2TAf7IC3DzwjZPuGKAAuJe9Yipo7XMLJRkC+iIVWaq
LIZcumGjP8ueg1q7Mh9rn4eKGdTWjJ7Rdexd5n3RRw6IE7cKpkIXYhEJDN9wLbEOpvx8R2SpgFwB
WZEPt3I6pupQzhZwlbiq6Me/T+TVOGyBxSkDU6uBAghApWNhWMF4W6DQEpf4Tza/nt+PEq95FlX7
2DnGBqHlodfW5/8cMhO8tL8I4WSNZ5XWwx6RIEd7yOiuoxf1FBZGtoTxIm1m/IywmZUYmu5u2MZg
x0neFxkGFjpxnxZ7EFc1i8VypTQm9BAXP1jsi114iXpSjkpUYk7k6A7VR/fGRrQyiVJ6WaziPT8w
cHS/cQ4t9SiAhfARX3zOHLWOh4WFfNRuY+rbavSOGNEqz/+4LdwtkhWJuOPXyQvLkNrtDASH3YMu
fRSxj34TxQYdGEUwql1gpAJy0u8kLFoIvBiDrw5FxyepDSgkCG5QS6zn8IeQ+ROGcaD7OpDQNx34
JQ0/RUInEYUM5kIzoMk0gq1+UqKch2nBPB+E4IWNlUV9Hy81v+Q+a9azguClYHqpJb6scfBCeayV
OOkyvWKMyeb/jC+KV8AqeaSCRNguW7Q4uFWf9eWu5/oGWMuaUoFCCPhwtkf/7NnOb02Ym5+2FKYj
zXRbj5h1stHBlkTupUwjuKdkh3VgVmIZ2jBtJuKtUpSxxA8YJc6N/13kYKXPElHP4LjNhPez/Ebr
uuBt2wjt9lsxREpDLgsoovnv4riWU9zKwoE6p+5yIU+1aC23WIj5tSU8zmxy4pHh8oEVnvicc/zG
yLpQId8vxXBuAsJpkFYBmiv12cwkssYp0XrN7KGNIxnOuBXfSkzwroBcVsGGoUCwbmrc69hANqyg
Nve2Tx0y3IOa0S757NZniTSj0D4Azed4mE+RQWYVJH6AEyGDcBiKfDegr4xIsWV81uOEXjPKNQFK
bnBaLWfledy1S9j2SQ6yA0xWFdIJeZmNDHotcttmg0EOS2djp67nQJsGRGOU60l/hdTD+9RVdtW9
lgdMQkBi53V9pO4H9R2/vNPgnIbwerQzM6UkQI9qXxEM2xcT9M2K6b/v8znbqPaQwAQO1C+JGJI0
7DXswn+Qg96Q+vKilRXD3QfnUJC+0ID7QZtD1RVwowMeMX6zTRYze+OSbP7QZNHSilIOCfUzIsq8
n6lzcLk04AoH0LzMhEoUE2fFjq7vU3DgqYXnYLEtwyQjWg2SXNxBW8MHj+F2XHZ1Zu/e/SXiDU/b
o8hg5yiFw076XeyHHBrW95oTYOIZjPnR6hlbEsQq+mLqs7UeFDha1pQDzS4L544H+INPuSFsYDmp
SxPM06ZegCjGblU8UJEchI/IJbSJeOb/gRESqeFIef+I9sA2+7rjUuiXpfVYqLUUfdGm0WsjsmfX
MNSUXDaeTR5WqNw9ajcTM2bFpQ/faZwaPHBZPI+vMmA01p6a8nYgg3iXHzqTRoLgDdgU2hZecMaY
f2u0e2L3C46ISQi7x5Kx0e7zeF2ikoApvic2rSLYNP5YbqO7reQNHthrFadNXBt1Ls8bzv1yXEnQ
SF6bTuTGVb7qIFjCnkVvrnMlw7omRNdoWrEtvmwlw1OmChTD4pdjPMe97YznIh0abJnQeqK8MzZ0
IBSnU+DA6kvUMW1ZoQuHiHSK1sKNbQ9lxSq3tHmsScUP0AAR6zDzJt0IzXvnjoD49YUWkAlvsi+j
ba/TvXVA19gu9+yQoMkwLrwnEL7OvMF+5r8PC8rWQk8WirhdFyNyC4vkEKGqFJkiuFK41LzK7TlR
D8ntUQ5GxMAQq/V2zzx6Hc3q7Zzi0zDNGT+DPWMin9AxK/rBaJBBEelP7x/R6cI1hHuOUkb5RRql
Ug3uuFhwu6be2n0NsQK+FeMS3g4cup8+GG9THaMAeNZBb+L91oEXyIuE/sniKStcHRhaL5zGJTNF
t5nnw7TIPNKe3rVzCpfvh7KFfHRreyraCP+RDgn0gTPrveuB+GV/VG2+qp2zJND++5g4H8SpWt1b
rrMbSoNI4Zij5DL63qqOaSOOKsf0SWZotD3xuhJ2+IY+w8nlS4Cyk8x/fuJa8yl98T70yCzeM3NW
YpSY4L1YNUdDW7qEbGD9csbLmIa0IWf8V9/n/iXOl3iyNFtdMxriLR9duK2rewWb4zM1ogc9ssBU
yJHHdcGCURiwmyMg5s5EPPPX/baIevAxZtzPrXqP4JGIxyQq3OJ6rIMc3eMNe2wPwsqjsj1MVWv4
G/F3EP8VS4v5eiXMfDp4mDVqu5LSKJ2kc8INLCMTfEX5CswwF9EZgpb7rDPD3KXhiX9XyTEQ08Jq
yIfWpJk5IZZpx5IU06oAXvdQNXtyUpE7JmoSdC8WLc6OuAfKgXZoRC0dEG9sLDAZngk08Y6PVxHN
03FE42gHYdF+Sx+8jtiahvVP1lo2qGN28Qc+D/V191eVPfEYrjTXniLWLohiHLcdRhNOaG29ODtP
n6qeOPgtAW/uA+/pamr31F3IBgo2s1L3XPqp2zp8uB4cLWWPkgphYnMkzMH7w6ouxnd2mgf45bnx
FP6ky1xBocGBj3ZKfvtVRY0TJwDFRr6ONNEgKpA/HauOZwlBMyYiW5cl7120uzgKBH5xKZW6YIiQ
c31vfzVF6ygYF8c2TooNJfbHiMWhQ8z+mfRx3k5uy+UEFOtVmhznSEer0DwWeVRoTg1vt4l1feHh
Jq4R1p+mbPH94N4YCxBvtL7ISAmcTmXvl6Isml5IwNj1BqeNuDWhWWGs68nsEJ3SrVaTHs4KKVVs
n7QjJ7nk8XB3BwMjFaseF6nz7B68JOAtOnVyErH9tAgcbTwOZ8EgPiPsuaOqMN1yXAz2qejj3jfv
GA52DHylIwd3ZMhPJJoCXMG6qlDLJ5xWPMU9AHTvz6FcYZyhBRxbuBv5wyZ0hKxy3dqsZKznF4xD
fCNTo1iPTnS0z4FcwD+A+S+eMeQPv3hqKSvD+rhV5ERnPrw4fDKoQKpeZD3d3iKQA9/KKEFz+gwH
mDFhlDwfyAtLQaVOav+cuKjmut92Lc4p+Bj0a2JAerGrJr8JglTLku+8rhesLH9Y2i/WqsMDKayK
vYlBSFj+qS4iLow8cNZSvFcuLhqdPCfKwfB/6mp6HExJAq2ALb85jkWkVADPrlaa5OUPLOo+1622
Ee75E/h98hdBy9ythrdtkrdaNK1qdANgYnhGqTKKEkoooA88BYSNfd4T+jn+4b9OSgXrf42lie+D
bBPY5SepxtcwdGV2NNfktg1SlVZyW72tbybvM01kLCdK+q+qWz/5eEHOSqJODx0G+HcxB0spNsXu
BbpXO0BTZladwUvDaXGHlgWayzxhL4V7FgaZ++Iupsu3DqbbHeZ8O2ajsHFEf5KpJswa4K35WQdt
bX67Kihra1BkgWATK3ByaNOD2X5MZpypr9/WXo7jlmgTo6Y53Rag9zcYejum+bInwswhxdhmnv3u
nx6gWLmvG2h9ErmtnDIm4J2xL4+vLaBGsk8fNF3Hca2ND5WSt+qLg9ql8Ypbt6zdk+FEBQvqFECg
pdFcRZEpZj9PRZ7P1QlHckZ5XtvwuIC0Z3NIIKiCALvv2Xd9EJoktZKpuZ7Wvwll4NANWzYdnld8
R0LeOC2IQPTIsQIOimBK5LK4wzz1Al8WH0Ym9IOzbtAT4oSGdqm5hGbYvq0kU1ATXP/8lFdYwJku
q5d3UKCNt2ietIRPQSaTzB3Y97MBoAJul1qcVFdPTk3pGkq3uGwxr+kttDdopIqnf1rF31lzHJo0
htygP9NJl2sYOQYzEFgOEl9fu9Jwy/JeRefotEr46b6PnywUHB5uoICbHCpuWC9PC/mH4QB3CcPp
nvPHOUe09RlHSTCUuH2YhBF3GsnkL5896PAZBqd/s1gdQpE8RDI4NTdp8pyLtEiw0BsbzsMvF8jl
zpVGQpnCj1Hnafai8Xflm/kpO3XVvyqIoBSBRPnhxEZ8FV6MvrdLO/MgiljW+eCcYHg8pq0+dqfb
SSkVIha1PTZmSeuPiSDtO2lz0wLLEZz9wyWGknBwngI01Fde/ecdgvF8+s7JUB5JVnSFbJJ8zdzc
JnPnOW0LiMiJQ/4XV4Xdk8jIdGmO+V/M1C5QT6HfRqcyb7KZ+dyIEKPnsEgIquezEXIEHCQX7f29
yoPHKxIWEnwZyFy3xWyeVAIg4bksEDB50TER4OlIj1OwZp7gHGocPQsHF9+VJbK5s+8JrTMrN1CR
RCJBJYLbvIj2KX9463WnnhpxmzuWOj4cMfdS5XWwYni2g/jeP7FpirWHsq5ZWCxzJufBAvu9L0wn
PqZfVYPWwHDYkUqIigPtTaU+53Ai0s9ru7VT/cBDSlxiqrpmJ1zzIl9cAdI9M/O/iOVDNhmdb+y6
UPxAOvNMVa16aWuoN9rUTwICZNXXJnGElf6BzJbSsdw/TBcteB6bWyX4oeYBmebQBMJvInHF4zyf
/hRYfE5yF6/uvbeCFFRJZIYEzyCO/PhkTXROEcIOjv1GJ+pLkdPW6V0/dW7KwLpAjQsmCpilOL67
grqTuGzs1FKWoJaxN43+W+ejGXA3mLdbjdMXWWoRJu87udDJxt98LNHsnz+g/hDMWe2j21I7s+SA
/sJMiyqSHCK3/XtNpqd+Ojzr5YCxisAmkhY3RW3OYFA3PbaJRCu+watI4X0HlCTIJoTo/5dr++wZ
XSH0zHHzpOy7O2A20y8TfFRCi5s4CaNW+UEwQRtBkX3EIs65ebmU9eQOtgxM8YmsQtU2vwOAHigl
npzyr48I0r/2MJ+MN9LImExRU3CasckhNJ3AvWX4oiizizUlPx/9rgLnxEP6IJZkDuQt8XV2YeZS
L42vmSnsXlQw+dLt4FVOU9sMz4kPCP547ZE+9mR8e+AzdaKiVm9sBQF2ZvrLZydYDgC/Mn7B+TyL
anJQ3QD2inYTwj/vomOApDG9AMpNqwIcm3ArunUw0+JUE6UOb1dH1YB17T81YnS6n+WE3h24HQYi
8hyKSSjfiEbXAWcPc4LJJPs82f2cZjZCnZD1UDYDSDRKHA3ofFbxqzXHHgcA9hIg7whI3Vech8Us
RRQLAgtQ1y1VTxC5HCvvWXJDc+E1epaX0Rg3HKdO5fovNwWTfqfJ+AjEiexP9YnAKD4VXR5LGB20
WU275Xd0CuHbid38rHFGlVenJ2xLdhPU1c0XG3c1Go+NMJ8c0vC+8SoDysnfzrZOim0u1QXyhsIP
tCICHrIDfix8g88wrQWBZST+Tk0+DzST4Pw16KzPhxgVIqjZdTD80nIi0VuabICDBW5D0vaLcNbB
eKS6JYskw13UsLR256CdUlz2hY32OyHsbvCxJ8hg4HUjUL2HvCEg+9WqMcyedbdz177UA59ctVgq
1OCX05rMH35wGADoFVyidjkdZXypETW3fUJOD91PEfoyekusbuFWYL10QTtxZ1FiWKDADfyFXsKt
bJiesN1B4ymYUCGei2/KeNDo42mbDAeShFuiIGmyVz0djnXs8ZNY1NIs5eeI2sQuneviKrehLWmb
U7Kt2U7BLwXjRtc7AnwZUEkF1p80d82kCXbUi6AyMEqNvc1kmIad3S8I2m8BJKH2JXZNrXY2NpdX
Ichnsn3F5FQZXz/Y1sRDM0YpLDxAlHhAyRMXHVaGJJauLau167G3z7ucIsBFhM51eVEA2Wh1pFLI
OmQt1DXnShqSHQJpy/Z00RqVVEoGX1Kl+SeIVcqa0wTUiUwP9spA53ZGBZcCMtn04IOCu80ZjoOu
JGzkcSMErqocZkRxWyDPpfXULTJFsJ3IlnUTFmx+VpxGCWTcjT0ZlItcMYxcxhAnS6VNP2lqr+0g
2hx//pklk7f40mPdRViL79s6HoCz/W86ObhXva2zC0SPdgDCwNrXWnOM7Eul/rzRGcplYHvNhb5a
KH511nn/Kenv03tt01HOP8242Gn7LwXNEbqYD9pLrbqtQIoOiYsg426CU9wWPr4ragIFSeywRyu+
InoGO0wG1SUBEOGxA67SvXlwg44Qbkt1znBjH20/c2oGlCsmEot3eM+9e1eS40Jwo7P2BuoY9+XX
ej23oHwkMzyAmwzoNkxhP9+6RWC0bchhI3B8avpxL9TZkcnBqZ90autTB6XxIAf6xaNKIl5GG1uz
FyKYpqz48hLXVDsSL/ElVwmu6clAFrPb93GM+fIFMkUdz935ovkEPV4P1/87qrsKsKCJ7XIgIXwi
/x57vok/Q/eEOTlfVP+Ukk9GXpjS0cGL7sqQv6GcP5SkyHexBFDbqtlSjHRBXOPnoQU1dl3rd6Ea
eoIM2LIbQm/2WfRzxcPD1H6vyAWktN3xrxOYFEjCvFr7G6Go0Cc8IgsEGVOtLEAEZWGlY+HSPRc2
jqPEbD1/cREAC9kQWPIeOAsS4Ix5cXfs3wWaNHFnHQ3xakLi7HuwhfDIS+3ziUsHR7QFm5IX9dHw
Sij+tVXui6GSAJRrkn5iw0og5OShjuqQPe27RArdnzOXo3cyMVkA9AyaanezAaH96tbK33/Rsr2y
vMwHEgDBqve+UamCHJb3bgC0UjuObyvRFd3AEIYrL63ftGRGcp5zJjgRUj73RSe8td6hcupCVmE2
U2O8jOO9AxomClzY/adJOuORDpiLfsQY1x6qOYrPMRa/1rOQrXgFTRkoCWjYIxg1KwNAdMkREa61
Gyn4BMq3hgOQtWIwRY/aXwvDFiNVIcdrC3IvZRPAvrje4Vr/zn48QNfDuk8TgYrCUSyQq1BG0wrM
yrn4b8HN/Of/pJMvfm83ZdxIqeCxGMtSWbD2pLXyPRYUejaePv+t+XyWwfhFirSP+HcoqUsLqmla
6Wk+w2wVnmEqdH6yRopiEqA0to9I8L8GJxKsBcOPIHR2JEyHHIiDJgMRarDKmBx+weI0ngEJza9R
IQeX2BiovOqs+8JOv3tQn0TS6AMUzn54XzEM1kbRX5LoPqhU7a6i057N8NdTSZ/inlcivMfL4E7y
97+Cx35jpOrZ4ZeUHgbzwQuoLSPhSIE49zYS5JKcyqgb7/BaYsPlMa8f6nsPaW+0JlRVAvA1NDZh
967L6nQOZjyZNBnEkQcVjNfZYnOLR8YnvLFJYET3wGTTehU/6yu6Q7a1uTeXSNZZwJOZ4iOMv96E
MZ98TUdv3Q5zEO6rMqIcn9j6ohUYzHhYjhY5TQrBFmRUu3BHlo9WUtwK3PEa1vWIUSrp0C/40Yhs
ezi01Vx/xEbqIfteJcexF7br7AKloVp8SE/eLaPVQrs/KmvvyfVrgAfVLHic8r2apfVYLOvXExP0
+HdLNnrAqDCQ4GhTUyx7zVQBbfydS3fgvgK23iqy963hJNOhgP/umSvLo7CjT8kn6Hx73KPmAsRd
fZTX80Z5efRnhxbjIyC+zMJ+lU06efYEeLwaB5kv0PsLnKsP/S4butkZrBozMrMHWv6RoTW4cGeC
uFxKUwoBsx9r9ZjveUeFk3RwReRl7WSFl/QuTFzhqFzzj8OA9lRgWrSgf3YXjYtB2JCAJEwZ+X+P
bgxR0Oh1z2Xa2XKCoOdY0jL04fgE8cL1MvnNuv0971HJaD5Xy5X+xKl5wXeSeWe9v8qBtEas4ZV5
ndLFH5vGewiqxydKvCRwYqGg8gDLJPD3vTnXiFiPedgC7+9rJ/j+q5YjwhDWKsavztEBjNUwiB1Z
HyRHBto8IAk+XJS0QO0vAuUV6Tgiqhbg2n/O46q2Uhlhd0H7b5e9BVDwSRy9Lxs2aLELBey68DQf
UcxHeh+PuAQR/V9txOS9GDorrjCjbFMqyZ841y4Ym7BrepHY2KfDQX9NAKOHYXr4Bd24RZ5JmARK
fFJ/gedKKkvsiGFiOqNkjDIoPoBbIlXhSRzq9oOLBucQhhtXfDdWVaZvKA2MItogMDJdi6Wg7q07
22UbStVonSWvC5ywbrEU/JCjwXLtp0SM3rsSqT5Fh/yW2F6aeK9XO6UFxNIDkYcoQBwNOBuiq/uu
raPXQpYd4/tXbN2AzQl9L//CXo5Dmn3eEpC6FZWBV2a1ul9k6sP/u0vxUUyvk5BgrGahlvD0pQiD
hdmyjIkZ8xZP04X9/5m9kHbWvn2VOFkFU1DQsYjyiiKsEZGhKMBdQU03qw8KA+gZwbXAtJrGdV5r
zFLh1C1Q/ENPzIAALWpXcqsizip940j2erxMcViLganixb6N1MA6JdwTXgTFALE9Pl+WurqA/H2E
0iAWLiTRdOL4iEmERuw58QfStTfu2mS+itFOT3GjwtilxsgGVbB7HsBEVr4Ren+dYNtforucXnXM
ECVgvgQlliJlTDRMfTTrSrMpjZvNC07eVukBW52/n+ikgBE5Q5ABcsjmlJr2ECHlFGeGLSZJjxxi
m4WTOKXCLd+5TT0+K0ctuzk8GxNi9Bmbg+Lyr5cDhgcIT3awxPi7umdVlIASsvoTJdT5AxmRTBO9
QE4r8yO1WmWCArcpc+gLps3pq9kooe4a5zyl3LQMOqabZf183lNvu3sCWrrhh54x+56eEwopvgQy
de2L29NwIEpKhVXVsuqOvJ8aq9GSTojB6nxW9oLFL0J6/RcO4t7G76OkcQuRrYXEHwkdo83R0Xxl
UQkFFNGQEpjYAvHJtlBDhXe6SfL2nFUbswpCo/G6N+9iWS84g/4BH7/9FxqF42Yq9llYKLsj+iq4
jhS7KI5k4BfU8Zrm3xA9LsR8Gd6k4YDqSDwacos39nNxoADxamyIl4EK8JJ6zXDG66sZXS3C8NgJ
npvHWPqGit+03U3Ak0dF4/SSFsyx4+TveGVZLCtgn2kPnSupdUuLfPjCMnCHCJtzlCHwL4orocv0
oTp7JOoghoWFPkd8gi7RoUu7USWdMGld5f63CMsvLwgYESvgDnPoK+80sEfQ8328L4NKGf88m9g/
El1ZHXLXTJJ5z+KiSkkTKubCQWzpnpCOPBY4xKliYrQpzDmIuX8m+aXxuoqSGcMK1sebmqZGxo/a
WPZXMcgW7ECDvjd3tAylmAEqpaemuA0CqNAMRsZMvdnq/t7I83Yl2/Lfamt2m+7wc/SYnRGLKNw9
0HRMIyCF2IIIHLB5qWdTAn7ZY5mzakRYyy5b8rzxPMuJ+omR1ruyvTSSRUdITlgdTFgv5aVoAVuQ
0QFRNRIIWZ433g9en7y+D2OFjwr5zPydcL/e7yFbD/F2EYt9vIn0BN9ex6vDylQMaJlTZtAvC7WS
0j5gU+eofiRlFFDmSApYLHqdb2UIkU27Qrxywt89wNxXlgUwFvcdE+ygRscCF5YcZNRPWK4dulWc
cHIaWkM+/Hn6a5VSqHEL5ITwna7DHQ2p+/ExUG5FLIkYMGPkbri5tM7lDlwy+5smr/ZpMF94Yd7D
XSXibENUsk58D/Mjj+EGokpQLf2Q+Ry5cm8yWUCg/58g3kHBUjfKEy3QiU6zJiyrpMuwbz41yKzH
RZemPP/Tp3Ojf0NH7BaFlwwWv0OghYBTVS+RXyvNBMmPSj6cXTeZ5f7AzMllsarmQan7BQrRmrLN
nKD3aktIBVyX94tfB17mKxju/L9dWPoWmx+uMpmSq7nnYKiqdAHweS2atsGE7PhdG1TsWRJens2C
yJnE1+Bsk41cKdgSe5bwbbgGD7fbX/R9qYx0Zz6+BtpJA2ufU2FYZJDqdPJYvYeQX30SJQoMEZFP
98+YkMplULZjYlD70ZRMiOND8GPR46HHGdKRjhsbbIkqGU79zr4NCAv1u9UfcyKB1WGv4VMHlUdO
eyX5CuE0Wxo29x1iXnyp9PiEZ5OAPT13kjG3Td2Efxe3uAZLVZOAintQdZRBfLOjcg1GkWgl2l8e
LzrHUxUzdOkhtXymPMDyAuWVvDFt5bMCXpLPqlo0SnfQQ74az7fyQGGZjnGbsh+TXV1YkJCNK7CZ
Xz/xN/rjD7XvmFLCBCPHmiV3oI9/ESc3/YC7OMmEdg3UFTrp9/zcdjNF8A+QPr1dm6bgRwrq6Lxk
snokr2W6TbsofoTPD3/YJJHoeFm4p99nPRM0VPbRJnrIipnkIjav4mLo6uk6pw+lI1NA0lVA+LfA
DoU3OC8ex2ImLpXf87e+QWvo+OigKsZJl+KeTzY3hfx/mECkkdYq+YinwjwOAEgeKXjAtTZNet71
eN/qZwWwY1kgXNQxRzo9O1vuJotrh2VoMKKL3vkbnY5ozkj/fpHFqH0RUmH194HIEaIE6GNAC4Wh
fgjt/+brLeSZWc30C9OOFsGbytTIAT+n9XOzh59tBIQ61QiWzv3WJzIPd3JPl8he8UJSzKEpWrel
/uxlMwDo2EMCm5FcU/cvxZt9M9cuxut3M0EpvLeCMDKv/RWxi3RWlDBo3Wtq/0uct9hukudS4UKT
/XI55Fytf2WDQj7hGwmYp1dmSlHPl/qDQxO+W9TiWQ4YGdeBZ3mb5T7QATI9fput4dmYUUmWV3Ho
wHTLuit07olFvRlg8m/StlAhfjHAFXwLS0iQ1N5WYZQmQ5J35D4geQUBLRcv6VEQxAwnUkO47ny4
c6rmCLBfk/tEyxJOe90bQylaI0nR5dushyXaVB3S0txBP7X3HrhA4577nBH0n69QOfsEWaaDxcRQ
g/+jpRxn9pJdAAyfymiurptSQ8U8Mu2zrRU8cW5XM4UN+p4IEd/glMfU/FpH6JwwjDCyQ7EaEdi+
PyOPBn4j3i0lpPjUXAiHdnpNCR0SPcN72Mq71+xQP/OYpp2ZgOXgJxEzDtQztH9KSxDKZSDDKqhV
R2gK2bo71eeemieZ/pmq8ZB3ZsLC9SlI2BWrfq3/PH9o/rbKdF3BJ+O3aork0taI2z0wzCRdJTDI
I6mprVtkbsadY6JWwO5AqXXPpKFBUUA656+3O8YUmpErhAtRGjlJEZcp20O9zT3Oi/H4jIv7+xTo
6v4N7hOJF/WabirRFWpmVjR1HbejnmL2VTVB1qrSlCDm9tExCm0SY8YZUFSaHMvs3abakAeP5h5U
XS3BzJAKjeTzkZ3SVIXh94Rrb+HjXqSJiGy8TmjGPR+zzU9gZ3L/l8oHu6fdN5u7tQ1xuUNbFI2z
BFiYCdw+IV+yVqBi9uy4mgFw6GXaCebV5jQBsLu4PliJOD7haY/GI4QEH69Kkj1BqdHlEIJqIFif
yOF0HTGq77+QavT8hGbUNFWHCaSoOY4PRck9+Kf81Ud1eteLt6RAruS1UJrFFUjBxtksTy0aYo8a
BTYvzQJ2uNEQ5H1OylU0jHgJs7/O0+ecdozndqgz4DU7sEABnoX9bUa9U+NzuDQB+kwOtQWArA8f
7YHijzNdiIqwF3VfNU4fwborKIz6k/ifE1Q01YCroqOAiK0dNNvOdGvdXb7RLSkuXV4dSaAhOVmT
1XR4WhbqWsxIL945/ewhKagIN1DzVR1uttB5yR+eGIDb5EpBBCUnww6HbwokyCk3jPqXYvRX1NES
HX9OlDXYfkdWZiJWxlfJOpBDG6eH3tSEoXlx4uw///jZ0/ckh8AmcMh/Bn2d2ysx9A0reDn/duZ3
ZA9i62vVNyylaOiTrmcXuXZUho35lgmPr0dgYFfoQOh+lCLGwL/UqR6SVjk6eICSUJDGPZZ5zFse
gvfq4kl4w1uQ2rt0P5DU4UWn7Ijj47MhAONN/TgDti9h4POkKKrojlAExI+um98W9K9V4dKRXyKo
ar/UYacaq5un8RmTB1mpBPPM/TeXwqFKhtbANDU8jHysUXx44LlBeMCWsqWVl13e37PLBoK0YBUc
Sf2u2z2RhNVh8BbZXKOjW9SqglPkp1KUzYnUUIydVVq/OqdQ/EQ6BuC8syArqRhGvXonyZplxW6F
i2Oaov3ATzfPOUoEgBgKjSl+3ViSCnBQsP15rhm+luEy9J0BCmB9mPxyY1Vv1zfPWKpFc/IyWVDK
NfaHwVYV9DSnvBDLW9Z+fuUXe+wgeKGS3AjNRX9Eghsuxd0yR/NfYGTfG7N6ZFymzPp/PElmKtw+
j1lWg29vAX6JJiVQUGe6HjApQ/rcNabhaq+HiKVcSqEOLMS/AzvShH5eN/9AOpPiS65wVICecnvL
YvY7/qCKb/QXCr/5mJ6C1Evwn6nN+PnIKOKz7JR2XH8J1QbJppn2DlbA8tCiz5qKMHXgYE0S88re
PYBhCujzvD6V0+kqwIsvg4EdYveFJBX6qhnUeNSgYpNaz7nNCoebLDnCLPkZhEvoPnM+DTR1BckJ
DEQuMOWBoR1zvX+QpCi0Cb2Epb/ZW02L1Ua3LE8RZKeIPMcUH62JT0eAP7hwzd36UuiAOSSzgzWo
xlfjm1mlnyRbcVp1Nm0BuPOp547DoVRwcO0JjM9bsslC5UHhRK8R1SW8qFLQHu0OzRmQ7BREuIdp
89+VHBB2yg0+sQNbjz88qaTHNi07XuNrSEm5bCUNKInJRSNSE6dTGfrrNOCRtNX5+hrHGVRqMkah
uTcuLQ0XMQyIf3kC5SOjI/Ayv0mfScMFLNVtHo7Ll+3iauZQ1Lf3Ed70qBJmq4pR+A42baurbO6/
EFIYiXL7SLiTQyVYV+4M6XNi/lQqPOd9hWbEGJAaA7MjmaKPh7ZNRl8fDZSaDg19KIXUngL7vz5d
mob879ETb4xW4jmqj7LzIIgtJQhwf0lLHfvXYeV9A27mX8z/RAtbAULqpj0c7n0L/4ceJs+ELSgl
DhTvZnTTEk/FOyEohz/JbeKBLbkyD14jjRWY83BGfatO633Mwo6dMIH5lvxUS6kHK+lXixGQk21h
hC4bpcFIQWR0Vph/NA7lSJpOo35GsIqEKYM1x36fQ2MD/0qNMKT+KUJqPnKfExSYyO1UrCTUFAlb
1ps2vlsVWcq8FzgJpKnisD8axS1SI7M9uQ/iZmfz2y8OuBPlY/IFOyXIkxvUDyi2F9lN4Zlyf+He
eYe7sVQ0cRyuBKFPHQljDjxdqCeqAN7w9GAT7SvH+sefDU2NSiD4xh2QlyWTX/8Q+RJY9Rm34gzi
pKIYYplnXhOe0FLwli/PHfJfVh8pfxkoc7vwPANH5v/M6LhkUVTYV+9Bj2b98jlLYtRgmhdnIn53
B8tioXVu3qHayuf8Ow07gSFcyIlt20WVbRxFo17S0E1QnKPNfr1oUn17ejieqkmaVP+FYzfOoKoj
VommxsR3MkVO4hBVGDnUhNQG/Kh1UeoYfi3joRAdXG/Ech6iuXzeZYI4FrPRD6OnJcu79+REf25/
XKd5GGimeI7Jy5vbeh4htmLBTlBT7wf4cq3ZjGobgD7TddO2KH0mueyrJDdpcoVXrvBAf1rOcOyw
KqgqDKlw1Fi6Ienr4bejMKseYaKKjhWTigH19vgbecDttBypVijb0Ab6mKnIOJTbMGMBnj2SbOY2
TUG7555aC0frP0yVd7S1RpJUWccXy1aQnl7z3KVaVnp7S41xgzdcaOPKwBY3Mckskbw4fLs54Yep
kYQJSM9g/Tpm9AggTHD95n1GIvAEzuCIJpw4qwcAgCrxe7mETagkdnnZRUgJ7qNYy5uwVe+JXs5Y
X3DwQ2199gm14ehf9oN1FgzfllTVv0LIREd/SNEB2yJ+sRiBumYZ23POQXsWraunPqftqtkcXwua
Tlx+GJd5dFDm/uHTBj1KYuzPbTGhpFlzeMEqm4/J09NN000VPFzhbjKT6iXN3/Zt2faNNA3W2c0M
NoEWPXLixvAelmvYlJSP8ozW4NvrJpi1u7SP9LkVNW481MNE0+LshM2IobvpSbS2RXc9T2CnjIJx
hGSIbRiiwmLCVQ7KgwmdvVdCCrNzbPWOQ54Dno58TV75wH+bAQLEWObJlzEg5ed5C1cVj3ewPpJF
teR+jUIU+j+pmF/ntNi/yVH/NutNW/CMcFSJ/a+vLEszScvQ+i67NK5yANSfj84XSaA6TLbn+deC
l82HFFzaF96kEn4+dYqZ1zd9+eLj/8/yK4Oty+x00WtvJ2fs/cEQMe2XVAJBd+aKLgX+VpvjcTyk
b6OmL8I8bKpzRQnZJBVqQl7FCjVp3q1msi/B49BP2dsU1w25GoHN1mAiDwOnnL5JjsYXdnyG9SBE
qBjxyKWFjAGk1kpTTUyRscd8rYeTvn3J4yOPs5P0Ke36RH+L6pBK8PSOUYQQf3DEnzOqFgcwM2Nv
m2yKtzMe6jaK5Jlav43UfGPDUMT9cnZ0iqWPSAqhHKkWf0JFDVA74eGVs+89V7JCaAUurPf/peKX
tZnERMsKxtuzlTVEEHpd1Smsuo1IN5SD3KepXjXPr9U99zGsb/cU0V7QcPsLrgV1h9QHG0GzFTCk
o+QLY3bz95jk3Y8XSicawDog7s7z/u3O6jMBPOEX8+mu9jEVuUy6KAmD2PUkYE9NElFVyIEJfO+I
Xc+8nrKTr/pVg57iQdX7q4yf+dpBQGkQYSMab8uettzV2CC66vt3Ajr613/eGc6nv5JDBywG05rR
M2YqSx+hneqLJO7ZPDfo5bMslyjYx9S4Oxa9fY1/tCgOKQr1IaOlfcOeymY1IMfnnoZyN1l0usXb
pHSkRf1rdBCnAjJGTx7330g19rWSgmflrWv1VPllHnWOlYNT6z7g1jhX6j/FgmkTsgnj+xMmV0m4
HIFQidoejrEGlF2pA84pNmGphGOfvSCPlu7icuuTigKKJAifjEM+ShEB7QmgyWqQklkyJdjLdgLC
DFoRGIEbjD8hDuUIGdvdxMfViHn/9lS5BGQASAAtva+e3WGWNGEEBM/oZCdQTh2pLED7sRXSUqyJ
pfwd6/xbQyakpiBA7P8C2AIBQzZ5N5RAlpyrA27OF8/Ve4z8hr0cS9lggtZhqtQ3XJnz3V1Pz7DW
+1qO2ZBzw0M85B8oBs7avxec1K5o+QcOWmlUaMqfqlXK/xDmkI0tZPaQ4bNSC8BOb5dLrhZ5Nz0q
dA2yUCAb0OPfDtRPKTHyElVMUrYX9ClmI9hPx2olf8kKu+H/OcHcQsO+2VdE0HRRo0IRXE55ReZf
KSj42LCVCBrT/MXY2724DqvSY0ioimH8gmq4O8VYDEr9Wekdy3FG45THFQ4C1djV5mWYK97J3Wxo
ZVkX0LSYaIWrHJUA62r2Ii1nw1liY7pDboygyOzi3E3ba8UA/XoPg6wno5oZNKW6UCI87M/LNiIm
ixtMtkvIMWUGdEDRef+6wTJUoH19vGj8GudHCdZTTlvJvZHtBqyNngWvMXtaqYU8aLTxXigmuIQo
oLJmw6lZ3BFfdF4AWJA0p46gSqUkNp8czhEF6v32eGfaIXKEz5Xeqq8GhtygiyrYVWdKfAIbC38d
n7vayjzBC3w4Ijrdk4MHIAcwD2CaEddkoqJkgXEPLvrS7pf9Xyg7SjBF+WKfqDSWNiWIdk7Qr95V
/LLrqUFs0vi9qwhdQXXYJm+o7pkL7nNdKPe0RINCjVKJeun4SrX7InNiXoHqctUiT2RghbTIBXtp
wYS3FvMiwR1VQjntj6/a845XcKHZmcd7AtcJQRteDFAXJtj/ADiHbZZLcSJH5gQMLGpuCBKLb034
qpWb+4mtsizDTmpyA45CnnA384Letu6+H89RKCe96gSXHzWHbfCNDA6AQ7fPcWyGkmKmCckMdwcx
X8Y4uArd5XgKrBddy+UvtpdBf1WX1M1aByYH/g9E6T0oyDwTe5wC0ric+vXRXlJGWEn2jZjuoGBF
au4vI7FB4bCmuEg+8m/RE8gqKCoGlcRvmoS2jUhlhqv4LtoCl4dMAP14i7aEvSiQO55nUNILaFVY
VCP3xlOMT3hyAC7tKCxvY8jfT5qXziJ7/nAJAxdwUbSkFUvZCTHKxJ/khkTfqWDD1LO5X61TvU+i
fF3sLydguV0hjFOts8S0QyQYWH65YRz6rtQRuspeZCq9PwYV4/HfSgXXvIzyK35/WVKrNVuOuu9p
/8uPl9IF5esK+8yHlMc54ckgNIVPcjR0unTi9V30+EuwIVR4NIA0Zk43CxeQ6+/ZFViI0ftpCztt
IbxzB+e3par7If+yzru4RQSCVCQbfVakAMM/Z8W8e8FpPYp60UWvXR4s7e9b01iV5B1KjLkwqNzt
UiBFuA1qh0mKfSleWjTvzfmJsauQmMYgaftJJ+LUy5Hzjf82qpIgAmauV0l83DiGyazK8pKVdqKo
R9PcuS8/QCQr7beoOMGNUhtvStDtKaBSD3JFLLl1HOHYn+bBSGGyFBfNwuKXgRniRCXfFatonI/v
AEGwivvxSKvMkxAZDJaWlDyKxwJ3OyTBpyf1vxAkumcwdNEX2VcLurkJRZnp9xTPCIz2mzcJ8wQ/
qE1s8xLl9mar/9sw4+pGFBP6XYrAPEo6AWb8d+xaBQp+4VIYmqhrb57paQ+f/YqaqHqu008thqwR
risP/crsMAZkYFvimpm/8MpkFyXM0iMNmjAW7PBM9/QkMXzjvlSKcjDWikvgaM0ok3N4G+e69xc7
H81mqygGjMFSP1n5i8pyAK8oOBjc17OKbnOY3LKOaC3FLoP5oxf5gNFEwyvOJ+DVpwY5J4Ud8MXG
WHOt/do4Hc5gGbOeo2Mt/l9cl3NZ+YngNfgcrvYsRPXj5dJwHymwHk8Aqj6G+AN8UmobgXnlwELu
EBtEfI8uchES4oIM/P13uc1p2I4vcmok1goDGU6yzRdQliMjG1J2c5yO5GOnvzt9Xr27yO45AP10
2zuUDSSVV74Vt0bkvbDrbMnGqAUZ4omvrdj8xj0tq6MOxQzNazal+daAkYlgqA7Br7uU6yIRQtoY
ugI9agHZEM8O9sqfQpDbaFc2DlCqgR78drOdZ/blO0J6demodw1rCbh5yZqOxdO8npUN6zlT3oeh
WtPuTJYOlgNVNchqwjjM/6QUSSKzS77AtuMCv9i4syvJAJlp1tSUNjbExDiTpGkGltDxDPit/bTh
lWg9yf13tBNU65XaxY34S0Q+OvRf1m+w/wsRIeQbW3wEoFvPus0AGO0a2WeHJrVBFTHAZFE6s7Hi
OwGZC9UGVmbOK/vbs/ogbBGWiVd8yEvjuBk0eDcbPqNK4UY+GKQkRp1w3aHs8TU6qfJ0afXdCPQ4
m/t2lvCJm5AzkUAi/8upQr6x3wtag6dqvV1jKsnQwIh6YQYxsrIAYr9dUybgK6dwoSPx/DhskUkX
+Wit3LX2y7qU/VR3GMayIkl0EGCJ0QrM5e8zAG5WrVFa/v/2PupedOWms5amlzzfZPvozVixO7Xh
ih7UgFeLFhzYalRJ6iErfBRBqB+RTWXhAcjNtqM0is3d4V/s9O/oUxbCNz04SDf7BOxka4fQ47pI
41K9y5vxJCfxcQ8pQpM2zFWBaJMviEo0e7ODKym+xfVAq6oo2H+Cr9L5wRfhICbca+qTuineQv/M
AodUNzbIY97T9169tP6OL2wxP4kEAOzwA6AGYGg3GP+I+pMdmOkbReogp/Z6ZDK6NdnM3HBZi4NZ
6QBY4P4oRWM6evdmMmxzXtRTXV8oxJO+D6Ndl+dCVE+biwGju8PcQaTfGAelpiVQFM9jmjge3njv
iaDIz3DOyLcQd+X7mhA6eiYA2oqiycyZ9zE96UEbLYs6ua2tWKYd1uA1j7vkDj7Heo2J4v0c8CbY
xmdXH8CGdkS2OlR+yC2ecmGQacZkAdAvWxNAUQ500yXVE/tCjt9wvVsohuahXUCI1Xd9S9Ukw1UA
iDgxppPBjRxpn9j7jKw157u6m/3HXdk6Wm9CBBRF9EF0aPyzk69QrvAGu8bi/UzMnflWk02HDWnB
IA/TjzVt9ngsvDHOS0xycVW9EjWNRHPwl5yQz1VK/ID1954/D5/aNfVAb8Dlfcd2TbDaRT55ef1A
82tkwLUtxnjz37S0ScMZlAmEFScuGAA/Ysgnx+Lb7O+8Oa36sRcn/+CBTd+la8knNhgo20ddXZjf
qHHMmMOYHBzPmRS7OtUZYRE9WVgPgpCB7EMyvoTx/ZG+0s63RgXXyzkAUPdIwNfBmF6wAty/YgT5
1vAvSIukUod81qVGFFrQB0mexugUBwqvnTZWgHNtS8w3U4kDd0bXa5tAULORJ/ncYktLqgdf9Vae
zaYZDRxiFCCID43I6XnuAhuGNJBEK7juBQ6aMjeL+Irp7+NXfCNaVUFcBxh5YuZGpjCu1iTuF2zm
fuZy6kKaMgGmYWwP/eBfaKUtTBLPbqkIHmnGu06LDFwLq9k9VpOdOajAkdB+H6AJcDNMNHFef3Kb
nhleizZJSoDwcG84La1LtHl1y/y0IfM/nGQ+RC7jocQLOO5pqUFFr5HHZTfbJixXcEcdCLIx0uq5
74yu7uOa/KhzGFe5MCUQxkvNAGkdrDRwcnJlzqdXTnwRGOpIwVltZfUSYXJ7WkTw7F36VoMEELcP
E2DdBjWS1MBRVMvi4KczVeeJ6O28aJ8fx2looozmBAoYP3jOjdyzEpqxCsZh9c3D6dTwuMgswlTo
RpZAo2uy6k1l7MGd2k4cQomZQcyHSBvcz3V/P6by3b9JoQ5WcRp+bE3ST8Kq5gUhMNs9YRaRXKss
ul2fnhvfk/CEzQi106Wu0Qm8CFWp0bIJmcLoV0u2LGiAuV28j0+0Jx1l3jDqR4m4Lj1xjOkIGDpS
tZGUyG5NPW7ACxDct4SQrQ5RcuehE/DuBpZYW6+F8lVlWdnXCda/v/uxvN0MqBZ3q/MxjYDCPg7B
1P6ivpzZ2wm42nnEnhcYYayHvaOV1V40N6ypLbLR1iiuZP2HQgNSUn33TemGtG1rii/6MZtS5glY
7VLNaxJZdOc682Ch5iuloec2k5lMR/tLNXwhYwd90b1YYcspUBi22jAmgRI4HHYQoDjZ6tuKS5bF
EE3HjKP3lAKRIanpg2gxAeHGcrQjwp4z9eNjrkRQvxaLCHH0uesYNJtoaWKaxpzfOXNIbfbmviQF
tHkfHEpkFBcdb7Mazno4lhJicL2ZDAQPa7p8LqGOjKEEz8xxDZm2NO/VHXHLPaYhL4HREKcWsvs+
q3Q9HsHFUeU4dE3h2tzE7sCqp+k9MXI7ytGBgztKxcAjuvnMQlPuT499adzfdPZfalPJw4pRLIzL
A/pAJboZFw9JqZ24ky6jAzU8xY7bltEuq4bWCCZpV9Mhw8o0vYx3dkGInsrOPbvku9spkKEAzAwT
YvW1xusFAcz1psCJTfvnlKOdJrEDqz+SB7cysj2hhUl7M8/Rt4KqefSGyYWkqeRAIDDYEiwfa6BH
z2FB2kj6SesJWzIEqN5FxMoe/+0l6LJ2K+fkAxM3RQ5XfgLHK3Ggh3Z8qDp3+KFRz2RTPG5ah2Zr
wIeaCClSuVCSW7VkIUv4H5yGypkPyrtYhXlq4JSkaZDAztloc+43jGYJmfG55F54G30ZfHItCanE
/Sv9zGjyE1gu9vkDYZQboq2gMCT1L7/Ggg6HbS3pwLt/vNDW6S5Az1ZJKViyxAB4g0EJMEWc/V3H
qqkObzMXPermXO9+JJg2hLFMKCnX+hVpsf5RBuO8gBL7XpdIwFhhkHlUMbaIfY4f5AI/cClm5V+f
ztunl8uqu5sBeQU6tK1u0aqpi5LrXPzp3OChyy02Aeswd3Jc47Xk5neiR41qe5ydt5w7AdiFCe26
98oVBLtTmzRsVOeYO2yLgUZZvPIBLSlYXM2QXQO/M2xBr9HLre/pozLjnlUDQpnY1CXYGgQBQHvl
NK0bJjwIQWbfFwxf+jdVg9TO7IH+wur09F50Rhy2T7krDLP1kMlFM08WtT6w8sVVMY8TJy6u16Hs
IRvc3xxmlZ9Y/LJwTuAzmnXifQxGBAEHSCPsTRWHXZSKPs9ZRjePX9HUD73OOnXRek2WcTbXdEET
jOW6RhhpieTbYmQCx0Em2dFH6HHTSe1au9tdSlJMsQycjOPmzqLQW2qWDO8lYgNlTe3ufwYTh8kD
0Civ6nSZYm1yLoajKfMo2T9RaxNybDAkrpUO7CwbFEIEKznHfyVz+lN+uH2pMa1J5gfaGTaJ+yeh
JrCNagQftU+5DguYWI5SgHPaCFfY8qM3Bjyhy/bwT1eLGURvlcRkUCBPIE+yCg6dZhnGbGXQQt9v
tJGWaAG0hFHCZrFnpwpwfMUpS15epNUuLBUVG1gvlvbVm6ekKMsDUrUEpfXgcVwFTAuF888L9H0+
bBNaB9b4DGenz5UV8BTHZM+DfGG1nP1soRHTxUWDeug/4XC3P8R/5WdYKP5fnEXRYN9xIJkWE8rU
wSXZfzuBQu+JgaQRHHBIpMuJtKA/qVEgUVTvgX5uGh5L5vlFi8TtvTou47RIqqJBvkR5xAH6uPWa
uiVcRYOEDNMC8czU4dIWqdmQtpCma+dJgtQOIRW66I4uy11HO//KW0m/ooUgzOhZ0ThOtYLR8LkT
LRz55kynUYk6JH1bY8m7IRzIiKx+Ny13pCaOPKLYujviFklhKuH+mdtSj/726lk/NjXK9o1TojHW
/otK7U3gZUPbfcGjnFX+CRLJSv7BVcwDktiJ5aHtHKA1VgsjIqmtQtbTwzjYKLFYnMwO0suHfbCw
eHsx3cmNF2CUs7atfUlod8TziAD0mtDYv7g9MENraMaW2iJY4vBEZTJxMpKI81n4qOesOeEolk6e
0RL4oAEOEDfVIoeC6XCecjNk/uaLsXa14SpJQAtSJTkEdR7zR8oKY6z41aRBaAbnQ6EnWzoD7aX+
1oVIHOoL8qso3lmZd3gL6SEM1GrwwQKgrDajO1cLt0rTkciZTWWBgHiRDA9+KbWGRbplFj8nb+a2
Ld1vZsq23yWx/esi/I26O5U+Fwq3roGUkKNXSlQoqZyOi8ytKXEEyQYqXsoD8cPngcu/F+zyIuZY
Xu6dFuj/GXTVssqKvMVvCIH8PUr2OA0Pk0BuiyjF+8nCTk9C/eGUqU9ZdXx4jpwZ7vGYarvGaxxE
qFvtOITR0qecW35fDTHDq1HvdissGfxB+uUkddQlqlDgRapZ1edWiFIo4tmGTKHvNZ5rfw7cbTgr
UnKzuhzXSawtHiwEreIG2cugUSXIMSfiVA7bpAT+BFbo65lCMjXwXn5ql1JTqgtziuC9hFekCu8z
O/CNfe+x19TTorZrplefH/5Fp3FroEbcz2L3w6VPCVjotQQpvTQSm139VneC42xUA8P7ERImaUkq
kQwhNoiwD4rILHpRUtPKgiOMWH2Af8uXgS92bMW0/hr0vlEGbkIO+EuF7d+OGCzOfvQdXiXOvgp4
GF+xcFqjct7tSPFTlhfFSc8z+JKg80Hojjec10V9a1TlF7KjDObJsOwXZUkAjWXWk/P0xcUcumyR
YAYN9K2GiIJUHx2SakxbtvRP8jaoab9uRR/mqXyEbkYhC7HTjIGyeLWEhBXsp8/2C7MUXJwqnZ8P
VwQXaFhF8hu+GIeIsNDnxfv015xJ5eTuBHMaaNsatWWXhgB4bie46YKRRggE7mSz/SJeXU1iF4JI
C/U1QHI/96+ztnEIy1MbW9n8Lg9BcjDWWpA9p2dv0KJofRtLj4iC05HrRnRioYDAFzrGV8LX0WL7
qm0TzRzKWVqJopv+DTlxBMvTEYBltXvfO83/MOJHX0zFEW9KETt5X3N/kN+ObJfQdnSoMdsdRUCH
6zVPmMLf3hjYlR/1vPuktMuKMESc97JtiGUfJKUsmeNlPQyhwwKRlPKNo28XobUzGth632N2ivkc
SnvZXTZ2CVOGl8GG3swBC65QGluRjBD6gXocZ/UEMrYtrIy3E50+WYhu+V0DuAQ8EsSV/ZzneRWr
MFDdhPTWYbPvI92qKhwJQ/7VOwB2yKILOTnox+NFAgI1mSUeC/G9r0LNkQd1ed7VgmRhyNYnWYk9
uN6jrZtOdjim8YQugdVHTS6ykXwYdBnFoyxKDCrKCWX8tLBp8h77WEUJks21Uf0Y6nmodDAq5+9j
XM5A1wS6nNGaWdtb4sTvtjOTFqw9ECuRp98u42Qj2nChVtFbmw7JO4v54FSzlYJfvk9hq2OTwCik
hz990GVNPxgCZfefMlymTxkZ5WH2rvibWMYHLANoGTbHuvqITTzhXEcZ2ivvYbiNfNiw+yaAPUka
fXx+QXkpSTaC9FjS1fu7AgVhUaCEaue5bK++9l0t98baHrV8mcshX/ny0LlFKs9+RB3xhjce+lDm
FGmLcqf2mj6UVrsCHic7pEJi7YpI+50INY3QEaRuyGoFa/79au55adbabCzF747HjelaA2iuQzDA
4gzSHISrAQ8Rnj2csdloDVqRp2JUnGN8KFoCgKlB5EyZx0v3ZWYUrWrx1SJ4F5rOopQ4Av8kq7xu
70hdiuTwNLmmlusFhuafOmiZ7HbxNknYSUaD5NUAxyODe2fN5zSIXcJ9Psb5W1i8r4WzkintRP5H
X/DS+3Ja/4OeYGNyWuXkq+pw8hldPh5+dzyOD0jsyNUcHMpTpxgCIaqgCY++R2DCuBQzoMEd/6N9
rebOYPajcEGxEWjszkxh1uPwtlYM9t8u1UGr65D0PBeGwwKZfchxIkGDVhdllwfoXpjFUD2vKYXN
VAuDLb0HGaCt9Cj3fgBGtKfVqOi7h6QSI7CGXNFjEdG/4UOHOhQMtLY/vfqPlH7HU1jipPhs080j
W+bn6ZaoFJqMS+uzZ+etk67DNXHz7ZPwUVtUDxgQdem8YxS9YISb1NEYQEyovIb8YZ9BkOtqp6r6
10n0jnkPYX8yCyk325JPzhhpi1aieecRNunHAj3a58WCF6rXZw6F7Bhx62TKJ/HUWbvL10Zaf0g5
fSxO57TvukfdE4wMAc5GdWrHkLXRzwYjQgtSteyQWfP4gQ65u1UV82nu/Kt9gtvqNHFNnKSUPBGw
9U2ik8Ho9vMkjGH0NLu/uro4Qt3CHKu6ExCYcyBpn9C4/dGSLnC+lMm9iPIZgOyS0lg5PZFsApKr
gvT49RCYN6iEFllkRgaH5lHNVNbp7NqqJ7lLKSHlHWKOh4v4nzhLltMXl9wPpsKFVH8JkHrTSg7T
lahFvwSazxkAvMkKAOdW9VMdlKlqQoxvbICmBKgz9RXFi4W5L5NfJQYfzmNpN5JMe47dLOn8eOT2
SCUTQNEyxbsNc5a4RBhJv9bTlp8lpRk2XJuIlCljAv7tlK0UAK2/bh1aNY4MK6sXySzDjyEx+Uy5
vim6wNlmwX264NlhkaVxqlEPtsLkt1VvT/DXBFqSAZdqM2yqtKhYOKqf+hAaV4ltQEGSiJFgX8AX
+ZF0lopQZ+5cJNvkx4k9j8dqAHworT/GDirqBAgCj5QouB4T39Xk9Ip/3VIZIvsmI/yhfblay6jC
fTVSfBShN20uCyJicKzdr4NAtLdOikccXa1la2fLxy2X5z23oiJd72Vyobjs08szaEbwBJaWe32j
0846LsLYwoWSqnHW9oqZTAbUiCq5encIuXB1eVXWEr1I1xhnykP1P3YeiJV5ajygbZBYKvLrEkLt
Kz6JiflSuWRs9cP7ViUlSWeqhQcupimMDFXE1olTEAVZ2Qx7+z4Z1VmsLZanXtMKgnW09BjwyOP/
ZFhcwUpSXk9SeCManbr4uvfQM6xlMoipGFnM9ezywciY8Dhd+IKB5KFEsDbMnttGkt5keHXxIFj0
dlRC/zR19kvh0pkiLhK1Tko3Cs8+BjGEFbakFoR3Mf7CV2knvXqZou6/biUOxzR7lpXX5Lpf28x6
64LbHgkzyB9m9PIVr/t8Mf5mz+I9D7MxPtV41QfZa62H2vUXQBzD6ZFhhxyuC4iuhZBdgHzd96VN
nBW0xN9EwfQsvax9ZvrcuFCwTZK01gbDcaQXKEmpy6WLGw0VyncudqG1MLAL25gcXyM1IuFkpDGR
8ifxeMaOm1uC0aly2O2oAkVtNO7lNtLXXfTXut2eHz7KITrvvvPdGgtG5lgGIaXQO2sNHv4We8ow
MTp57OnSyHhnE8UktPymPCoaSrCfHsDe14SXrnDBgdk+SO7+dxuMsulNiX3le4L9AFgYH9TyrhKM
i+0PyVyPZ30biTpp3WXYmXPRRKAkb1vG1b5lj7ZSQReu4ftyDMU1CjIZeJM37GAkG7rPXCJx+qNd
trIRjVI+Uwu8bYC5oTTZey4nTA7yn58KLp74q7fxv8OAGPzK4bVh+mGeRHOINyl/xMsdywzAgT5K
6UndMxYjUjRLuUWJJWHvnh0uqxrb9rTqGTLShLuXRV389S6IXZk92gC+XJ0GjAwXIY//9FcKnZHq
5SHgSv/2PaLjo1rhf7vRzguVjWXkdgkFx+bQeXOsCJjSR7Rb34xLLgK+ELu3hRdEC5RdPYE7C0XP
8XsVm3vwCZaMz/q+2RL/JrcP2xE47GdTveI4fRxVDn1mny1JBVrL4GVEMsBsNf4P9LpjD1a5Vkl4
ihHfB8PmjXURJfW5RhNR2qkpQbeKoakqF+qSWos2LnoKj4KxoHWnt0mE0yBhPyMx4pK3Q04hI47a
+oTqUap43dUOcRpmiMQjON++FPsxZqLUnUHscryA9peALksfFrvWg+egIstrRdIkdZJcb5I5boey
UDSFq03A/4LIBbiqrXFqTYZY1NoX3O4weVLIZvC1hCR0SqYsjPCsSVmuYHinrga9iXhv0dpEN1An
VOQyj0EKBrl6RzxCDoZCCtxVIdCzD+kJQWaHEpzQMuj0Mj39MDwKenG7rOfN7jJSO0mX4s89rK2r
TEGzbie1wqwwF4WuoH0QFUZZoGyKN7zs6Wpn47ZFYefnfXbmU8XKC1C4Q66FdOeFMqZvVI6HuJT4
sY+RX503hix9eENyAsGO0vYyzlmXV1aUc+Zc00V9HjDFz8jGR4qN7WQgadW2dGLESO5eP/HcB7Gh
iqBG2fKZ2EvrZy0bXZH7vUJ3/2UzdUAUQPP/0+dnImKsqs4Pd5yFVRhmImsttSWZoqovEM4VjIKC
xGE/hUaMaKFW+ww7Jb0CqCgCGfPOzvYF+FVovFUloVamN5TEC3Y7YNhzY0Z2yWk5FuEsCndaS0FP
Vr8Zg8/c0WW/XBboYUJf8/h3xlvOx1JdaYBVxLIrnT9eeJ3QKXcT2XBceY1cy2HmM4tiK/qcoB96
vz55BCFqiVvJWfts0EdDFOXR8Z6C2/9MuKOxZsTFM3jowGSyjK8DNfdlKLu3HuPvjuhmYgfXRD9g
ZHgraFSJfYrEDO2U+t0TA/PxEisrZYRVlC4jhFWPXxfF8AjhlvniGsWJDFm3dxAOLL7wmFr2Drzj
rV0M5rPTe/BKJcJ5MB307d0M3nsrP6SWFfXnN026RfDL3OAHsAofkTDTC50cyFRkS8N6G/cvjXEv
2Ru7eNx2SXSW3KGeKZR8htEbsXpSG4AcaPrv47KED4LF0AiPdgvmjLYLuqJEtbpysQkRAltCzVsm
ZP2d8QpiRGrXlgYBHD+Ql4B951j1GJdB5tAjRL5vsps8HXAc45HSAJphmMvAo8i7J5Mbn0lMnHEY
AY7Dz5zr27GySIjoV0UZP77Wh31PTr7mxpVSn+VbpkoA6CQZKEfrb0OpDuNF71ppDflo3yqF95Y9
Z+mpl9BFWrLjhWAJer/yxA9l7vjDO59SJ5N1yCYWtwDfQofUWmmi0A8vvyUR/dxWy6dmwBKLR01g
H8WOpnohpMrdGkns5lX7KR1Qx+Zltlk5pWMYoJhYq5FNEG0RPtpI22CLAjGQuVYNlXfjebe0ruFB
pBMTpWYOjzpKu/2hVKC8cVOj4FtfBWUKWL/fFZbxOWNqiQX21Nucob8n+NdwKZ04OziOa/eqdVsE
yKMLut9VCP6+fzRc2Z2Trs/4+T5oxfyDqKgVm0QO04AZ6JT0IgjK/6exAD3oJZpl0WKhGXbl1YtG
PcUc/nqhjVdkpR3Dre4Il7li2oy9h29IbD4HxKTLO5K2gbTrFLmRya1P+FeEqY1Asz9l4/kTBvJ1
ZrqK5PgnbCMyUml9+9gIp1ppUQMiJc3NnKlPSjQffgQ+y88TtfrGmlQpnMRcz2tIGhz3rAr1sOo7
kCzGHC2lmoWwKjyDqikSbt5eps+3xCaSvqc3rGSGroff1u8UoWQuTCnbzr+0Rgiiaj4Q+yJPTXNc
qdpIgymmZfuJkTLmXlTOOlPrUesjhxlQqHeogRpo2c8p2Njl6d7dacXvInQ6qWn9S8vhUepN6ukr
MKbcyWdNLKmHBcCOt7Yu9PhsmEhn3XifBB8yT4rzR9jz7B5cDYjthcoghoD17BCYJaLPW7o6XV4X
CdqdSX2AOSQG8I6gZgxH7GtU2TVUEbUqr55k+4tB3hL6Km9jYeud9hAbu7AGRtoR94x0ENocDkhw
M+iAFrAbpgIOrqIVuZ9+skWInmJfbzeUjAdZ8/4+VJnmgz35jQDOKbtsXajf2omErX6aQ50Bx2nt
TsYRYGzbijdchj7NWYZSn8oWm66moEl6dIg+M6R/WVTCavUmgxWYvOw1fNyQpFawsGQDbPn1rjcG
jCIMc/2Iud2jlkS/hK8Rqz3ShzyM5MnX6mEKTy/YtzE4UL3rLouTKt7S66y3K8wXWYEZ/KBk5TI3
wT2eN+3X5UCgSbdEJpA5mKhSjBah5G4KJmGaaWnMOwEDiVjQCCAcivjcQnwsDbqWfDzY37S83xzP
932aoPLlAwDgjNfHU51vky2ddIuPIxGdYJng0yeiW+0bUvHXeR+9rg2KLjTjUH/O6cMbDkUicq7m
PctbeYYPbR5lFHVXyQvQs2VuaVhaOP6oJKwze5RFI9w/g0rgf66ZT9v0AtCsXAHWLA7EIi2q4vbX
ObNLd+fdUHoSvc6Yc5tgvoPb1OMw+9cHJtJrYjusgh5lenjgBnaKGhqAVSta4TVhJ2F8kFgcIh36
iSeurhRPOLJS4WkDpx5SeYoNz2rmC4tCJBha/SBmaEkv2AM90W+F5JEJAtC8cE+zuZHzEhCyRLiy
cBDTA15Y5EVBFGSGx8P8lpoYboIo+j+VdGXlGtuM21cAq5eooogRVXLr8HSLXM+VXN9O5Use/aW1
dLTgHvEbrdiJ089i7OFDJPY52xrCthfvDI6j9/3KrDnyspuh/TLifTaxXkUSMCdZ24YJ5xrHjNia
b73wcnnqQgo1g9iGnHkuV344TeuJdAFeBa2Gdy5SZTOTSlmmFKeYmKI2MzlL2kGOWBswJqLd0f7A
uCzvQi0a7CInn48sF+4LB3XVIYapeITDzqxEUoCmRt+y/av/B6y2kZwBPm8XEdE8tPR/WpZmcBTg
cDTb6sDe6ypyfp2y2KlybthAu/FZaYS2PO9ld24uwlZwgbRPO0e0BZjtex45nmW5FGYqER/iwq30
4IPowGK6fS3rXGf6+CzDy17//B7O4R3oySXj7mf5lIX1aYvSgOpzp3LGLmbX5MPeibJGFieagAHQ
YWNYUgBxC+lFtnTeVzwhpYtdaYm1nppsfNDiYE8IB7JIc+tb3pJBqdDuG+LW6m7kXXOd02xfBHWs
L0V286Mz/kyFR59eMSNCoNE2jz++FYuLHmVHwujlzzNOprsBMfAN0nsHD7peLO5ef1wJt79D8Owr
KlriSJLiIMv+Z705+1h2NIRS7CJhGlS4OMCwzdljfhYgU2jN7UyWXwUHvT7HFXN5Sn5D1OvyHFi2
n1ZYlpnwEZpB/woGurR8dvSAVL9t05p77idowLDY0LublTJ3PUl+dErH4mhWFjrsJduBZL93oy9K
R1N41n19Na+uug2xEQWa6UWfiqSxTkJuufhQEyzJYyGrvnnMKf4nuLsUO+2Q7aMvVd5qXF/rT7aG
Yswkh9Ckm8jCXKI+SFQ2sJPF+dwpGjQmyEiGgmJeNOXZ56bnSd/5OEKid0tiOiF0Lp9u4XoDC4eX
ifyfrYZ8uHMTfyXV08DgV3lcA8HcCBuQtpJb8MCVI5D45zo2QPsFYv0letOl+dbu/CebMCJJHwP0
/75hOGReiWkYOOH5JoZs8KPye4oJfjW1x35EuFTYtB2Zlw5vBkPr409B3E6R0oYUwy/vuuvZy90s
Z6hJAQaZIJ7iDiSiB2vabK+TG5UP0EMQjd/bRSnTxfp7LOGs5XBSK2/fGOEjXifGDs6zBozd/C+Y
l7LA/4y9vqJnu2SagELuiLaNgvA0pEnmeyjoIvDjhsGgw92OgZlj0eZJi/qsIRIt3SPgnVSFGr4u
H3OU4O1R7zPbxg+9qxt1Kr8V9q88kvP0mXJgaoae68CHbRv3+6GCm/9pYdJe4BsoVmS50FMzy6U4
yDKPUk9gm9fF/tJcBddxz6wqzMR0CvW/WJqDYtD660Av8tSBfm6DuGrx6a1gEht1FQ6RVUgp9Gqu
pgjQ8wDRTNnFPLOMpegvApoLHcDIR/XMU/K4eKsCfo7ZNCFonibw73Tytq9C0kLy4FTcTkZsILT/
XeSFkmcVsw4ZYVi2tFpLDT1u/hcH8iAELgsLTHko3uOAz1b+VGUkjtptSyGsvYWYrhHMjOcrE4EV
68gzxf3CHjIHQbrIrOvk4PLDZ5rTCu0RgTSJqGNfJX+5xQws/1D+i4AIZmsO0WzqJJ8BrBNyOXEI
gXkLQ52sfzmFbg2wPIHmfu3NCMMz4YO2ohAnIM3L5OXwFwgGZDUnKr1e/ACamhr3z0cMTsT11oWl
orbdWEqOV8Dvx1I6sdyFp/4nn7srS/bvu7BZGN1VRZeW1B2sJjvvRW1zhMd7wygAn0RjofO9Ukxj
UlWWYVYUUjmJ7jJV/BOz2D0uFFx+MX4iyIQgF788byFuCRNevoSGXnke7nKbQiJewkBiMuZ6TKrG
qH7Bxs+HEWwNCpis0P3FG8W9mgXCGNz8yYyU0/37Y37iydgT/Zi6ZsIzEyMFEB5V4dS1grF1TuHd
q/sUWTszPYHdAfWY6qtexY9kU1wei4YBF2xtgcPoviI7rREpVi8i+Pi6di7PnUBYPO07ZkScerta
T7avZ2oCsv4jjYQ7smVdfR5B2o08OqmAgy6GtvSWFUeNbdFO4kezfdTjvFTdcBxvY451KSBIBqBY
KyP1uJEntiGliJPZIFoi9MQSOH0KG/7Ukz8ptL76OFmbwwDvwtHAlPW9DEGq6v/TkbBwrdoyQsZp
MfLgtWtw3n8JLm9AYFR9LC517nmSA5epO7extTrVlaoqMa5eDcjwu4amzXlAJQ4G+5oQC0cAFuI2
5dE5PHUkqus0s9uDajcA7SQyR/M9MioNa7wSJwQ/N+6NokS9y39fmRnWO7ZMeRYN6Xtw0wniqtsa
xxQmNcpK4OPp2MG6k2l+Y7wwsFRLfiecUnfVKXRdplqKcW30CBtKVxWKBtQm+2GVxrpE1vn9BFmm
s/z2DsW471JVJs9UHuYdBZ+jsUXwR+fWaA1HoEQhBEeKIRbc8rFc4QY0/+N4HFHkIuaetYfzMkFB
fPbMzrVbgljc1SjKMOLFOdE81yHJg0nGTuv/pw1dWu1bIelBcWZDLf6avBR2Jp15IN5mT9UABtaL
toB58zBGcUE+tYtvdAh+d7p77wuADY7+iqbJHVLS5xBCYE+NnOFVXOeur7LEHQdDlSWmQC0heztN
aRKpMr0D5Eb+8LOj4IYj+c2waddQw9ctr0S2zWw/6tQdTu7uD4OehRzL0ms0zj3WspnkjDvFyuUu
Bd7Tjf4ttLHyFNanC6VqNIvl7V3Lh1azR+ooZrbDAjOMY5Ay/pKRm60cHbJeyB/2/2lV8qGzlCz5
le+7uXroh7QfgVvpodnPUNfB9LvA1CG1jg1B0qlJcwC1rwrjjTTw5+t3rI++VAektd3Acoj1azh/
M3Zm8bziFpmmQBGMORBXmmnXLcNchw2a8DHIBI40dg1Y0ky82GHhEo2W/CtRrgqqmMI2RV+RYz3R
xlcry+ovuKXMvw+HHgKwZ/8Fmd+dJUg5G8zfKtBogyJxowPNz+wwgFMNey/fq5886vKMf8i2n/e/
6TpXQP/3SJ0ONHY8Lx2spg7VszVza/TAkYJcy63tB/cuw4kRObziacmoQSLWEbr72hZzORHO9AEO
u3IAe+4e7k5aBSgIvfcFCBnGT94EsLIzjfbHgWJ99/99DEUyX+nHj21juadfWeTef+PX+A4nXc4A
hAc3Lb49Xwz5YVCBTOtSnkykeQ1nTMAOeGsBnz0PX32ykAA94lpaowWeSXltxwsDuo3vAbQvwuGj
mJg9wXQ/42nITd8RNW/MokddfYsrdzZtpNYbqAHaOcbyT/nDCzM3EsMedCvkv4kMxthPQdx75jan
hCWHD+qKkTDm2wihDKST/MFNkexbgCr5sFqWwSqqwdgWm8/YA1q/CYDn1Q5zQJac3KOJMuYSxopk
yMJ/QsyAHg/xdbvXzFLCPfa8h1uHCOkt8BIQcbanp+xFvQEivPRNaZ4ehVwM0hdjsZKFX7tZ/+xT
2z1WN9zM8iZ3nYuwDzNrMBMV5ClG/F8Go3pUMPwiKjsjox+fqgrzo2VKKfuXnTedj1zp5p7SGKvs
kl1t+GB61W5gRN7ZmHepHbjV8Wf38B0d1gvgT4Wx6fllIeweox02QBwQ3+dRs4Fj9eilNDyYH6YD
BemjBVnllrB5Hd0iAF9NbHOjlQLpUTyA9485WyfY9n+JuvCV8pTlZUAlShVFLu7nM567MblOUk0I
AR+7Y5Rrq0wWOYzO1V1j5oPABTIzZcfp94Rg5AJsAiw9TfByYyAlxmal4Z9il6zp8o68Q4jKvz+V
Gtyom0gFCbYdm2KENO+x4k4HzcpAQo0Ws6i4NzoTBYO4TRegfTWgEjBeKqVAxvREW+8Jjbea3bgd
HypZqkWm2BdrUUWHeXJRAvBd+TQQPWosthCpltggyEJ5xkMI9bzUBDuGr7MC0IipgdYveKjdJLoR
eM2/BdDU5Y22i/vbrSyKv92ua6DIViKvoXtLfOP88vO5L/mNIJjo2OhBDQD1jlCTvm5ft2FAxyxD
SwCICfgEpafRXzzLCdgCX7kCdbn3aRAQ84ubh7T/GsaFmh0jM6+6VVG729DMIqEZIpnISVC0HuhF
mrqBh1Z45cKMW4vQosrDX+bWxDZy2ZaKJQlwfinGJM3Od+9oZbgINIguBDq4iFO1Svas31vtbjZ/
qFzX/bEu26qjHlXCECh/nM2MfpZppWdyQSWjxu16/wC9LD6x+R/Wgb/YJZev7D6ldgbk/1NP7VWX
jA4Ni0srdXzWoo/5U8tqFdT46LH4AXjFC4ljuZcMZVYUnxkVgBxwCAWfyFiDL8d8/1R9iK8gYR22
/12sfj5hiWgG+7Ufs4N9SlNDIxv6MpaQTwDHPJDvMbRGzjfnBLaosk/QI+Wp+qktk/qybI0pcdtg
IbQi5kDBK+d/JFN51EVE1FXUjbu+OwII8TY5TAsESHS3XOqHWfC1VNXChM8HHI+mJ6RGgtpigh05
v023q/WI/j7a8CMQnbFic4anHQ8ezzfbFpNr4nBoz0dJpI0uDhCucQhKBcnWRl7C0A7oBTDoyGiE
KEf2A/gvBjhnWPcgvE0rrjhdPrHYVQsu6qTjQDg//7zy6cqJPfjsdFVng7Ue9IcNsA1uSc3zFrxd
/+J/uDzeyxWYqqh5UovMCMWIXDdOftLpM5AyZm+C57bVq7wMev/fUtVfcZ7TXVk/H397l+tQyE0M
6Bi2SOqcylYuZ1zQIompc2RNqMBE1wLBuuygePZYCxqyRfaKZ3V0hjC0CeQwTsFw2hdjBz/ITq3Z
EotTyhLhxPPLCt+t9tLYzNvjVq06Z/MC+r+mbzABQLfovsYT694pR8oS75weOpju00CjAAkjiE7C
3bch6DYGIZq/K/Whj0KajUGvdbMiuaFqepX5Vc5t5kvgTiF9o5WyEs29TTUMttTW+r4mKv+dOWNn
BpjWO9motpqbzZNVODGGbJyhZ0NL1cH5CkuZt3UTVRkTkHPLlMkp81ol0+dwsUDIP396s80JmPht
dswRS4EOjUR0G+SDVM3WykkZhTsO6dfR/+p89R00uLrB3QQ7vOg38W3dxGjRrhXk8XjF1S4q+0bb
/L4qwxEEx7NXIllZ8Gtb3Hx1d2NtC2F+8poUuiN7eZ/+mxB7Cgfl3vGqHgzTcxsqr6qlXqUVR/M0
V7yLUPrYIC+VxTcoxUWrnLOv21DC80ItZnjkgdAptHxSTJYYkO+dSGK7ViS0OjMqic5CivvGddiV
3yAKfkivFs1K1/XZhpktsKjv61JEOMz+DR0sB+r6SeIWaoyRya9m1gJfbr0qsiLX5GiWrl1y6PzH
6pfIsKiUeuaFiDj4E5y+N0xarr6BJ2FBTXofQgK+4c5jSDCAS10vWTYzCmqRHGiFdHJi5A/pJimI
NKziFb2silDurP3oTZ+budgN4b/QOcQGV8Lc6q/DHQkGtI4poBALKp+LSTH7FD/d0w8bT0naguV7
Qx972nzeAttbWyW1RMkF6HmvxvTppDFYXtNH85EnGxQrGz3HQeBSS3tKksC2w11EtRdIQSauHgRV
QpE67SiZC2OdmJKgaDsPLs8JxaxEGHra5XoTfM7O/yANZW8W8zrMutdkOjuMgDe9WlUR9HkXvgEj
VdhJCjRj+5dn86NK+m5GjCzVWXuBU3QibRUAgwX1YhHNQkvFKZERbcSBKETXE7IYdJZFl6BoBLIM
/p+3Hjh6Iv7H28o8J48zv02STJI3MEqgj67qqkBBFw9nzBu7ZRYSqnkyEBaKhddwzdDfHr3N0737
8gSvY3jTTudDIXSlktRtcOkrMdUtCKXgbYo2wFe5hs8VEqySzb3ExDUCEa/Y4Q2S22NPGV3TVd+3
7LsGZ1rscQdPyk6k40UpbL3yBlyRhnLuRhphLSFVO9LqaV5w080PatgH6TstP66Tpcs2cbOdU/PM
9Zv+Qtzni797h8GY9csW5aiAUYLFyvu0UFnYsnjthJAmzbozR5Yq/4YGGPgxMh21GgmI6MuHC6iG
G4d468kkqTKxNq6j/T2aFEvHqomwMyHtXA9xNLn0QucPmKLkl0KQDC01R62o8EmjZa1VIW5RPBSu
Y3RYC/Lew1g1+vaBw9ij7xLpp5oKETJrM72wPzBRqWeK2mV/ojIXT0Sbbdp+N7/liux1l+1EKqh+
3oZqWflmowQjyhm+dEa8lYiFkZXasLCEwrXhuHEywlrHzfAifWOgZoPPG0rfgVF7lDlmJ1RvPhD5
Pr0RhEqAihRdamqugY874ivsNb8Avl4L48RRZnqITm24BTRHR9bgtdmhWdYGTTyYghlyB9jI0Wgq
xfuPnAiKv2rbrIhYI5kQhAqGk0K1IaJinIJhOOwMbm/9lhGPrqI1ODEIVpje5WkKptNrrnEpNHQQ
Lfz0JJk3V2BpS+xtCEOPv2T7bglp6SiZdvo9fudtfxu9w2AK0Ji+t3SNKhkQTWpiMG8h0IAbqTJc
XSBXoOhnlpqn/tRIpQvA2o+UpD3KkYiVdsfjUbCHmyibSZJUmX54lOZ6FM1W0ChNCUTqYhe/RAZN
9cMjdNaj05w6+W4a3jejRu7zrJRcFwYB1y6c+WiXzd1scReE4lwTER5DaReCSG92zNMTOVBfC4F2
4REmS98j7TBmxmYkxy9xy2ZUaRx2+DTR8dUgNDfMIBUULaJedYEMMdMdW3XMou7P+KMlezllBscT
OttQnXKK4rwnBK688+ToV8UqOA83OHhc6MU+gh2IPSzM7ED8z2A/ZCdpBzcNeDUefDcGruWyUnc4
r+nU8aiQU1ehqmwhUoImUYQPzkcfZEoj3QLr3UCKaoe47rhB+w6uaBtKR5qFbrrgKyCe7JbkyJce
12mmX/fq9RgYJ/2ug6VwFFLaI4HOvJuDuAaFLalcLSX1UglZWvP0GG15qD9MLklohSE57eaKp6z8
PNFFW+NzwtwR2CkAx2mO7aP7/lRUPWb3/Tb4OP9P8wRV5FNBrwhnzJXzdxKDj8qIojY6UMMqd7qF
POC1sLm6k+jyCqpMmiE4CLrcgRpb0TMm5qfC/gkCfOgzsVy6mpKNh33B1l/0hDoZOCmoylp188F+
lhNjL3wRiS/ZMS1gp3WcuWScL3S0AKUI6gMZn4cFchVpYQzgvzpPLdRbYNw22wuUZ5aY1+N4K7vl
vPlpkGCLJWH1V1oc8QWdyFfE2TzkQ1JsPjU7ZKO05rnJV6aq124CtYdaUXs10ltXXmou+ku9ZYkQ
9sI6ds0hs/IWSkmo1cGZolE85E4EDx2iFKwDqpDkWvTJ4UxiNsTw3MDm/aBKbLmodmr6Hr5h4XoJ
8XML8iCA3lh5HeE71IfOfvSfQNiGuwrYvsHlrhRJ4Ch6jIEU3D1zjfpPG4BMpSTDTY9Hw0f0tW2k
M62Cd65w8hciPi70djRaXFt6RCwpRqAHf4/tINbrdkU4/8SpYxetHh26m7dLRGFSS+mo4zw3qe7G
HAD5+B9VL/PI0yeL1Olzkp+YAxgWmulrfZtEapyD/izvCclK07sRC6KpNlqkKv7saVpo4HFyty8Z
tIAMajcsKIREfmu4NVjC+KrHjRmPLA50XJM/XW6MosjZWDHogMw/RN0WYicxCnVBemSedwkxMIIl
J7f+7OSn+7LLvaYnITQ+sVmp2RpQslauWFEAE6mmUiiKI/LhxOBV7PQ5Oi+EEW5E9C6ge9DO5URi
vPWcurKkP7EkjAf24wQB428XgNUT2PgCfmBvt9LDb1uueCBIoDT3uijSJlVQhmeIWnUwtGmPJY2a
sOkMKbMxJf2CuMNAjS0QHRUlAZVfLCU83x0fYl+iZboQGAfsZm+ELgqolZ4WrncX4V0wXFuiZ4ht
8AGEC+/mqTfJtUWEq4ohyXYFzwYsygyWfLEdX2HEfWgdi9OLisfd9Y6PPPAjS46fh4HyNksA+h2+
s/qlTO+Sfb4/Lfi4tFlEXvYjop/1Bl4RCNEJSlrPRMSS6nNddb+XvM0c969p3mkwwDlsO/Smi1eD
TpKCwxc480yhpQUDIgcvJmGKgbVr8PIoYrW0K3Ypn+G3nf54XVG3AXJLYqPttdyvC+7vYMpOXMFN
q5R2E7KF0+7VS/vf4B1eQPFJXuQbe6FGLFYOBNx8FNlxUapONRrRmqRqN6kg6IHsMzvousDEjYJl
VSCnmGyPxuygXz4Icd12REqa9IUlfzzm/gJVSKFjImqarZ6os2ZERvbsIphlUoi0ei+FVHHnjxVI
/JhF3MvfLX1eHEwRYSG8ArkFVSMzQsCjCX17MYqyf7IhOOw9cbKJl2la1Uqd4nep0PbCj82US31O
EcNsSAxRqBEAyzW0rBpGPGWFrlt/F0X8Yj8BixI/VYe048MBmTCx89mvtPca/frU8tOsy131aurN
bgpB+EQHam/xaJC3XwnGEjwqDcmw4eGfiYsBSh8ecq+EzCPYTITYyURM14OXVmhhi0v6/CimAe+J
GsrbLoZFw3p2g7rwnljeUsaBwQiIOs0PlSkbn4n3vonTN+/ipFoSvBDWPQEdq0eTEmK88scBvLYo
znbh7ZY51N7CThZLQiSLV2pNkvGmDaa7wUCAyAQv9M6epAEEidBDcLSBa52gUUb2dnzeL/xTNt2k
QvjGFoUE6gBv6eDSl2qVVvrhQ0yxLCijfy3K2n28BABkT2eQWZw5+9w11POacG3g2fgNFaUBY/Lk
YVRPr9WX98oBJrgbVH63iZqcXYCferkgTqg1qV6SZfvAXj7Ot/9st0D+Tjq9yD1jViQudfRi0htD
ifeTLw6Wh61yYq5wpCxJhRpnU1N6OMscSOPNloNmKMpsUu1iPBgj4Fs8RHAw7osspFDrJJclyvLI
XCBwXPxz4jrM1jBqbkPfx468yBIb1iNVCfE3rokcugrFYtH7HaMTuzLExo/xVzXPfTisG2XRe6SH
NTGodc2LgcBvmf8ZrIio4hvJbD26doE1aAriROLk6H5VsUu5ZnMAHae3E70yGZVilooVu2FMH7ck
vq0gVIi++xwrmAKfwLySSLql4U7YfiMCOh9NXGJKCogv/1ydStiMCw7Dj4IGKAji1mnwA+XSaJXc
nchP5da/UrPU/diXKluDbv4lkF8fHYHprzikE5RuEcnzWofyg0KSnNaFvhV2VVcF4NUEdNCQ2wup
YMMN9VYJg4Ma75/fT9oDv+WEThUc9YlfhxMkHWVuG+D6LOsOacpR6aoBM5/UbmhKdpP4hx4d21Mj
EczuvDSqMp8xB4CSFfuTvvZPCMwbEIdzV1WB8uz6cbRO1nU5C7Oyn8tZXXILNlrXZcxYGH31lgpg
1+UrBNLigBv61Z2KreAbpfRr917akIjbbHtx1mRlKPQ222RWJkIq8MYMu/L6HGw2X3STxKsESPx6
q3J8/G5cd1+6yMIF8LwAER3gZvIx0S90bW1DrfbXrbnq5DNjKJcAbXD9+FPqxmM25gtGWGQNyqE8
byEObn2ZXXXHlH9v25DEetN3m9D5Vcpo7MnhG6enN7vnTVAYNstv9g3+oNJ1qprUHZXp/zEZYwj8
cMcZKe1MPYyRfc3vrSY+CZEsvjivm3SW/ZEAuS8Aej8YgLw1q/DjHnYt96vRnBxkszxGcm/LB0w7
I6w2qUmaWWrmemPRSdKRreMr+r1ST5iRLsMhFTzmE0SDQT7NLYNOLLIek0h9HV0M1nw/BhLwfv91
yar4Rm3xgUSWu7//A/StuBQxPpmX6VzPY94WGNDwBkwncjudIYvrJmYkUd7PvJ0vX5DxUNvk55EY
4wrK7e3fbFXcc2pd/1dM+htcM399RNtQeqsCDBFdiWDzz00D3dea57D13YjBQpnUvRdS6YbC44pI
wCZiXfUWhGq2DBWN2hc5286beaeqAU6uvL61cDe3vGxv/2T6xzXGPz8eSkmHunq0TTgLt3MJKTLe
uiwXmLVPxc1NfZHnxwwIWCIIIgc/9zUy8aGeT7SnWIxlv0kEVKIHMRWDoDc7lI7I87amcCLR5qJk
z6X//CvBSiA5n/8PHQ78aFeRTpmDJPN8NwMp02NamiZigGweMTPSXsWRziA40dZ24ym7Obj161MN
Q9qxu98ZlLCnJwpaPWneoCCCJsx3CY16uNKspPTZTGg79YgNmaqdf4vkFqPD04bkkhQz04yfmgJk
92tkGVniJnaRLJPsP6dcMMtDW5y5MJuZqfPSD5Xu+vQX7vBrKOfQAq2rtnzyJqWqnRqgtighefFW
HVhiV1LbNSZOeVtLS5aUGQJsBmwryhd+QlVXS/Geg5lv9056LehMqth8F5Q5ODkVP+bnDqu7AaNT
Q6DHSEASBewRwwb0CXwBXv2Sl4srigu9DuGBToaVSsMSW51myHBccDM+APidvhXJwXy7E06BW+w2
+X89wNcqNzjwY5hkcmhymwA8hZLRQ68rNmffD3O7Nza6l9WOcuZIoqAlpdHsQdvWG+QXAPC7Br1h
t5l0Q9AzkvY2u0F6b/VwbNAkDy7eGnp6/6LM3K/UxVIxfEFfZ9zQmXgF9Vv5B/jPip83z+tRir5r
sYzzOdw4HfpdQ+p9Mm+mUZ9WxIUG8cACY1zPdIrWjaPkTaLEfRLd9bKuQpDcFqGlYvtlblmnlpZI
BCRPv4L4FebGHoD/TaMMjWEObZ0KCcu6MuMiIVk8arY2Jgv3F1IuY88rs50QVH0VL8aRhZB8VE1N
Vdkg/hyRz/JX8flb0qnBV/vi5y2QpT5uuCvsWIjiK3BFhD0NaZ+scFKoWYxCeAm/4K++Yq8eRev1
HMFz1lQbUuPz7bKw2B51Ak429ufJBaWkiG9ymFfrmeR5Ycxum7WpuGfadQ93sFvC7NFHk9DA8omN
HMId05fEPCojwrFIx/DUedu2JbXm4kbz+SBK5CepmqOsocFgQy7qYFh1PBFlLfnJYsIQb/Dx92od
cMfCvXqjwNOeqIqFOP0/FmRsiOUjf9XEaY4+ccVSJ37a6uYHd1mMcVc1dM2nvd83zYHP47VZi5gI
XpsHPb3GRcqkq1xkjPA1niEc2Zkp9U+OWR6pmNgs8YVxVbWkEkE6IxoqXN199IR+ExXGCzXKUFbD
8JeATbulCJ4pr51JImFuqclJiC56UG7xMovLOLGZ9vVLtzx/9tO8xu4jj10geV/caUIXJxy/cYX4
pge7o+glvGdZdzQhWrQoRhBQdVtlhRlJX3agPTarIm2m/5DpezP89WLIGRjH2YMu/flbHX7/wVK+
gG2YITBo30pi0lxASV5sqmNPXSRD/dy7lYlvrr3rBLjMrg3bBMNj1frUWmF0rZt02E+Z0o0IlSVS
L+iN6W2BDwWZ88R57ZtNOpDP2xFCqt7IyxME/o9tYvxdaeX+otJ9RLsw7oSVaS9H3dxeI8eDWlNC
QcqJ6TY4UeUCm51OqapzlmQMjpIcQbu9+fVAx5ftdWZf250BmBr2H0OXZZoMzx/BqY3Djb8QmchO
xITt4k4UytC0Ys/EUkBkEfnA9YNc2XJBl2zF2dEW22ibPYdzOGzq+mA5VBtIAzEOHJCppmbp5hxa
hezE+JndOMPLEtlcpX/9f/fF+AplZKhARtQHm4M2/hyaacDXUkaQ2cjfPQGAPHhAowGtKaUJHwiN
i/tQsn4dScAnnUqZUWt+N/ePItcBDDBY8x1UoQZn20xVr7GSbG9zIJL2ZhYApfdvmOYDgbvy/BvU
VXMecgrS/eYMn+9sL3bqs5BG8oLM+rGJfog18B6sHoxWZxERyKRvK0wsGbyLS606SwMiU2tbBXgI
DsAijnYviLbGhfltrcTKKHx+oV1rCqQEDEzvKjxn6a0l3YXLZQKTs664KiwS9wW9UEZJgjyNj3Yf
KHY2NdQ4cPlW8YtG8NFJ98Biis51qsla1rQDCYNLu914SwahyUmWz3FXCf9YT+h5mWWD2HWHKD7I
eL43I+AQy9twAbFVqPsDm9t6DY/OSwscBWVM1KQd7CNUW6rFufbVUvuKbawl5rxJO0JDns0ZQktM
/rIcqgXdSFylUwLbp8hpa8g1pCLB7wLBl+6bas+oxY3v4Jzil/83E+EwF7aQ4vfhTj7/Nd/GHvgx
yzb/wqLP2dmMVJx5BfRI3CZsEwZ5l4kXI/52RWMwRlFEm9w88ho6MeI9ESPnQFFeXh3Va/aOJ2/X
k3o2oPCVDRvWZdbeRbywIUx5gUrIVceWsAYYOjYtMJtMbl+8wzcer51zuOZ/AvR3QTnyLGyzTH2F
tE68MDzHv9Z+8/JANffRCn8w6DVKbwLo/gh2fBFkqSck3fwAUimMmCc9d5GqNCA6XdNwuFVISq4n
6c57tGgZdbOpsLFHwyRvFF/KfzgGhqCKxbnYNZZxMzlRFVuEsj/VyYH8P47/YJDQS9vf5GMj5ZcL
zz0syVtLbFoO1T3mc461AJSz9ZXW3iE21Rm7akOwSPc0NJRhqP79m4agjJ4E09Z6mG4mLwvydLiS
621SZ2/lFDGDuEESTwAPhJ99S9/4GrYDkts7EPYqhaCvCQgMCS/QvAzoeRmao3g1HHO0MFyaltn3
T+Rp9UQmRHdeMQ4sPqjS96UaDxhRuZXb9BmFV9oOo05A7Z15FqfYE7frbkALYp6BNN5d8HdU244b
cX+LauoANfQiYJdhv+XsftwCpHB0Y9tyy/s0RtTX3YkEszeQZQwR1K9az9bgg6hLcYJqhQ0TK8Uc
UjKjNnpqblUf9orC59PSa8z9ooHSkncLEwZCRdpzz5k6ndVLmlw7VPvn7XIxKLONyA2EtrqDAAyg
kDLVel8ksuCBYHi4ss4sjXC0wNsvH04sx7CxM7T6YN74pr7dXW0b8+y1fKksya3flQqGXeO7jbpw
53xjWIxZnaeXPKT4ugDrR7+1wv9jXexBio2n/sEBw7M+b6ksyMGLp3DlwB4gPw5tiHWxKaj1VbAm
m3OA4UOv+P4aJkEUNoUHxWea3OIizsFBkkUwVf8qJC+NadHEduv32dacSVm0zhzeL8MKu8dW++R8
bURECS7rPG21RXDQTtPPQt0Mhr8q2fuLohm7KmXHAvWD5ertYqW+Luue3pccoNVXXtOAL0o9q2ER
9o3c8GqCxA1+IfoRohD+sX/KhGXh3kqQDUu74r+j3ruRKvjoXZef6tIAw310V+r9ScTE2FvQudyI
wf08XGa44pQl8vnNBjgZLrAlXLljITJlYp/L7omuDOCKKg8zWUv4X9+7Zb8sqb61atkDi2Rf4uRD
m+AV4s/GWuqcYzQxtHb9R3WcU0pXSaESmTSEPGnfIUNWXB6S/ZOkh9vfKIdXc9udo0aIkkNXDU2s
KKo2eyR7TKGGIZJakOYQCWX7QLpKAhDVkoSWmrh+usvEzcPjtLP0DgWNLBVJ+5ayd/OUn5JfcIwj
TLvl7MoLhbnLjJ4lCK8v5GkCeI3ltmps2qVROT8ER4RnFnF3m9h7LYVdIHVddpuHCk0VOZ7ir94H
FL4rTJwhKAUz41h92JRQ1XiyVpT6p5gjROjUYoufknmn+u6/w9ZIvt2yvNiFMr1vAJMw/wvC5ndN
kwaeLkLbjrvrPWQ21wBVPgI+zhEqs0CpBJ6eQGoJW8+D37ZCNAgJ2QEw05pvEtX4Ft8Rz1JTkD1p
7ynR8emibR7JDLmzTuFkvvZtQtB3itnb593A3Rag8iEEkEbZVL7zoIMn7KoKNUUw8KGbwyDGbZAX
m6rGJvtRmzwVEPK33spPAtt6jAQ9a2fvWnbPDHoH2yfCp/ShjPH+6BGCDly1y7Vf4E+dpf7FzcLz
veElM3hB25+KhMSS5BoLFh/ngtFo2IFVhu7HINtcAhzC1NpK2M6B7yiUT0TQRwMDii0AaVfowHdy
+tQ7Vd5wMoqCJThrM18iElzzsCVnNFj4osdiGpRqbhDaLdE2jpeBS70qh+jlOpiLpK5GcxKpgn/R
GCSCCpeRfDA9V+OHc29qL8w33+QtMsbvViSVZmAr3kOkkzdJdSFJ8iSuy4cgG93t1EI41m0jvVUk
rtnt6zqMZrE8fnIKxBNq723LG0XebgATNtakC/03NrdwHHSr1no2h0Yd/10iy+kb7gnnJAvhThOI
3T3AnktgZyuFhembJem++sJTbDLFcjmFFxNe3uVXUciJ9J0dgRFdrGBYedpruMarEjOjUKPnGEtU
ktCBhema2nw0uNx6WvfiqlB08JRkdS9QmbeDwNOg7RxImVfTcmO8TIbV3tnd8wJ7wQw1qzyAIiy+
c8VLMFP/3Ap4hwVeXxVe+5+WlIZX4ii5Oh2AYpmnCeb0pQ5ppSS7aRgmBvsVTQRJdD+DJFYP7t56
GDaxeVgEbmqmeXVNUdtPOb5jUMnuMqyZ9qvXnaESX51yFdZfyELPwXTGf4V1K+f9osbdyxZf5B5A
h9xcmL7VGeng8O/+zTnY8q78tl+Pj2iHjJ2orHUdj3Poh0LEGElgKteFNvHIUbbzr2wSDwEyAiO7
yb9TUNkC2LTxTvzZ9ont+4JxmyNzkPUx8DbUZspEDi4hk3YpCYM9xK/hLPpcha/TNSsfKXw+SXej
qOnf0zoNh5H7q3pFBHzYI7EruSAt7LdGlu9MDHg5l9BNtQ31szfk7Wh4Mb+7r+Vvs5qFJay+uSSS
nejTZyBFEk+RP+Mfz9e3G+GOLkykCP1wbpCIzjR7eQHVlKzSeW/OvxyEMo3sTm1Q2x6hbXYg/fS5
GFZbFxAKKEnZ0G8g7TGAeA29RRlNIpo+8uSdbmREPe5pwjdZavK3GmXjzjH6gV2KBH4iZsQ9cmJo
eguT2Iv85OO/7O9lWJUDTit+fob6WQ4N9vY9e04PZgwnXBlAmlCLIR9Gu4DnCDJ7aIVZSyGZ7nrV
3DlgyJbV9aVx9AO9q0NQlwUZutY3RpeaNEHz61RPj8qhNNSsqVhJJO8XRlQcgrNMNJXTW29pVC7d
e249saZIM1+iUSemC6R6/fJpHrzfAM/zYG+k0HisbYvxRDR5QZWQXrbJpQpIbCkj9eNpGDh3EiIq
fbqRy/rCpYatReCQMCewhjE72OhJ8aPKPDv8Ox92pcCLZYtjw1cFHCyfWJPtIjYscdDwIDDDvTdo
NKlrDwhHgHKZEcAV2Cit99PZ0fn7hqoFqnPpnTQwiDDIwTJLEIGz1TPDDK3kSFu8DuE/DvPXu0Yo
Gq4JtuNFr45LnQnDhcDzraOA1fu0NCvwPZDU4KPpVRnJ1joUbyrgtqmYlzjjBX/v447itM9IqxmY
H67GwfoViWYjjT2Q9o7Vt8GQDf0L+22MuB8cYUj5NBVhRYZwqEiZrc2NtIIeYTXl7+X9k929S9X7
xIAjEDegh3dJKgjmNWhSoonY4g14Hd63bmIMhvPEdr+Y8RNR409SqC8QdDJs1XGUn5PIntvGjULu
dCywAQBstgHRltsOLAEqQ2W5ggIgLuG2ttEh9/xjehcYc/VXtx41L0Hr55N/IWfoU1akrTlDhbxW
om0LO1H4ldGzDIXBblNMAn2zfxZy8/U+oEIqrH3w2k7rxXXDB/UkrSunrbzGkSV6qEMiBee3NN+u
oZxeISusZzFEEjYl3uJjhcYCJrTIr8TvZvlgIUWNil5I3X6LATdfOMkTWGWr/uJ6+VCowpR8cUaY
LiZBUgaznGnlHmCZa+GmyolwC/+1f631ZgcU2ng+i2K/3SKl+4qm7RJnxjZnRqmY3iHyBJM1cU3v
yCTjwE9vErJ2MvU7PteTQAVdnRVLuXabEVX+Xixkf6Rjz4n9HPYVjaQFt460n2f7qredO6FrFMrF
tUDBPnpzwlyL3reb6YUJv8mNmtHScmxBVQRQw6h/HG2H1FQ/T5FFlmCsYl0JCJpLucaVOUpHN8ku
r16iZdAMxw6Tuu2aWtxEwxz3EvBRYJRU8wlwtNL0942KVkZnR/nEbqMnEqwzyUSkYN1HAFYuOkEW
zAR13OVUdW/8dLMUVcW83PXlTNEs0vioGrwQU6xgMjCTSRuoFjmhT3E5JQyjIU1Z2vWopH+Oz7gt
heVAC9Qr2sfTXOwkuCpiGopBBsbAeM6NRIOySXdtwxT6QeJ5VYRCw7go7w/NV39koOPW4WZ6J5XX
/8mHCYuJ5xXZTysOxb2tOGz4j3wVCNP9BBv3tL/cuKZNTgJ2slgEDD/BpAwo0GY+mFpddrC23bQD
Z/viHwVUuBaspyTsOgGZO8AX9hHSI35ojAPnVLQsJkDa4Bu40pCS3SrIPYeRbWheRB9VcJlp/gxi
OtjinyjqRPIV0dreGnXze28NdB3oiZ5/kLIK66/I4WLfZZ1Jl6n8Bv2y92L/3ypfuPLPV2Ml+VnG
EUj2rXgnxlselTZEsl9pOnSBSFEioQMwVeJDDY0XE9qqVD7IL73ItPzA/5Y9dol/bpeVLQhZvHL9
5WUjnfy5kNdh9wJXKyHTvWUif7yuXhugtR5fHWOW44zzwOfMNDN94OAZMCEngp2FTV4KA+jA5PJn
7yWTzHyFrHbxVSK+tPlMKTBg6C2xUksYMJl22eID3ISyL9Gbofh5NtheZOLc2VMTt/C9ud3TDxrb
Av2GFDqRSwZs4rrhME8uNf7wd7pPd5TKL2T4/YbwoarcV4BDw2SMQAop5JJCsXyphMOGEDWzO8Rj
GObJWdO19xI/ovwHYADQ4y4whOBurryNlUVF92e/bgL+it8+zIFXR03TWyGeK1L7yMm3gp8yEmyF
t6ibRBO+qFbC6pC2BxdGnLHqNFQ5+r5xWzKiq30dnQRYU8WAkmlnEJvvDwQFTo5AG99rJtzryQb7
K8RJ0RSH7LVzw6N4wdZeHbTemuCBr70GXvceBN8u6pmeJie8ANcjjOipJWGEoOG72bT3olQJdWNI
U8Jd4VBtoO+pE/bD0cNhUTpK+RgW33BazYzADwz17jNXlxhghopiCAmfME+2F+iL/bDge8YoU+qV
2zAoWr/3zCgElEKUXxi3r3D1H6W5Fq6Fd73fkbN7rPV/tO8z1UATRs4WZ8Nbi5J516LbqCz0IUfI
Al7hT190evqtyVLfQZYiQPkj8oIQCAQTVbkT4bJC08VzzKQ0A0UCktWirzLyterSEknHhM04oWgY
UCfabk8rGHS2oP7W8SJfRN7tsPDUSuSF5hubK4fhnra1gTbwBsxvt04KpsmbNQiOxD10Cuo2GdBq
9Qc/pmFgnxUdV+yDTRo0u1lmLqoZGlmerZs54jnL9e2SKfQuqTdkgaHDJv2jcjuk9imbHvCq9Pkx
3X91clOF8kmHPzee2+OyLHkgA/QFoyXkRtkNyM78MZhqDMI6OArH6k8O4hFrq99XA7qjYQ640x3i
KCsMJMWUmIPhAuJWeguV1+UF5zGBtIrEQVf+Zlg0chyT/KLVH2VdMRO5KjKAKpxDhcMjFGj8584e
gQDCc5oBBikgTk92f2FRyg5d7YX8j2ocQ+QeNTVHkULPbiK+yizev4iklrKH1zEsFz2yfKxg9gWW
XtEvYe8n5AjNF53qD4VWARkpXPNRLJhgb9Tinc0qJx98Xt2FKAa7IOVlRkG+y1YYbvHqe2uMhID4
tCHxB9xXJzTY29uEHi+4ULHNAE6IkQyYLlvlqndGTtnqZsHPK8NH7xPci4MsG3lbs/wy+VyLaN3A
mJ9yZRzbuBkluDJXemW6+vDeOPqdn3MXC8cspcaZCv6aWwbnXHpOyQJS0maGkruFA3zFcyCIQnzV
gH0txSqkbT5BL5uK5l7vw4NOrifE2BckHSZv+QWQy9/qYD73HH08gCYoaCJixZjITEZgcToHCl4X
his9DvG/wzN1/+5Q6uTCghqPIc0164esGYEJ4iU8Dm38mD2Jcq1ASHH1OyV9mxzsNrtjG8XiEN+Y
gEB9Dy8ePov6EYVEqYOLnZ8vdZeH0UetXwPC8cf50FFT7VxtZW1EAj3T8ByO8Y/gp/W0AOmJg0zd
PLH6lElQx0sXgBF236ikub8DiO4bduvSS2YrlF6TfVZZjnpv8CD8ocTUC9ZpmHSZkuX4N3pTAkjs
4XmUzsbMb2JSl5se1g8nG1VpZ5yM5z18lfnqdzioL4ZMSx3+YBZQAhyXpYjnxmUQS+N9bENgmk8n
5GPxe6v5/YuP/iYwZx92sWZjcOgGdkIPxxhR4+TA9Mma4TxkPokelIr8PEGthIV3FvGZr+4tIwA+
gzNlKe1OVJMlqyQ6a0h3fbdUDR+OaFlxnsE/yjUAZSNqFlw9FlW3xruFl8p0WEnqWfAN4gIM2S9I
nCyDpVmXSh6XUyKf9w4nhmOEGbh92TfFdHqvFRxlKanDW4Fw8NyNsH4BiVXyWxza9NLYYvtpJvWV
f0kBs9TdSZh6gFgDFPinIveW3WkYLs3Xjr+buOC3T+iWkO3YoLTtTSpIfIo5QVriWJpwA1OY1Qdi
JxN5davN9L2z2fdMjXVVFhvJ1csQ0N4IuUP8kGhqOVYRxJxbficRTpbs3HyQ6WLWyT15PmDERCAf
SOVWHtEBmMXQvXmTrwienp7PdPyLsMBlIqcGRUZdpgWuGyS5DGbEIceJuHa6U8g3oWcI9qXgO7FA
eBUcr6JPyRZfN57aDA3x5O8v9tSAO6p3zaXdtXUreAoWw8LradTPLDMB/Aw0AlJhSZWGKziLtvzD
dzBukli7HZSu8auNFy/JxsxKZS1S9WFfHn3CPYwgQeW2n1xdEP7yi5P5CPi6Fz7bybhwfKX7HzyD
aSmy02ny3tpnPV/X6FbeO7o8YOxJ8ovFcmpxFINPJDJajJX39dsZl0lhbFedQdvMgn5B5oi7E15E
ewjkLLTecW9hlRoTp7G7LytWIM9oCnDKSZQEs6U1xcyQ3VJqXH98Vnuq4vU2z9ozx9ttB/Vj8Cko
2f8wF8K0I02P8MkyyYT+ZZNWcOqygNSZcmFQlwj30geAHGbUH3Tz7vGEICzJL9bU6W0N2d8QEQ3w
eEchswZWqreGQ23jUAPqaG7xMGxLS6ifV0SU4diWlM4j7INJ4rfabiCgoW+X0tGEPEfJzVqdm6bB
bUnPJSjwvfd9aROvveXDbJFd/lZeCK0uhulUsIITF1EAe3Og7aQEAPF6i2MviC3FqBYSPKhMZhQv
msdHjuN+Jp2ehOQ5qIn0PsdVLz07WkQ7OwSTBqtVqqhA1KzxZABZ+QB0qol28em7KcvrCCNNO+7r
+c2H5hSjB3LiaHnnyhEsrrwcf96Ms2BNkJ0nZIiaqgfAkd31bYxLaQ8AaZ6KRtRlwjnl24M1+6G6
Dd3H54pWbtnpcz8Ff3bCiTHAb0xrV/ut0ztERz3DYQYrGPuIAHsa2oCY96LTvC2DJVOLo7gdUOsT
1k9Pw9j7Rl8/cjdRl91UoYJjbxEr5/3n/KabSSCPhTA6h2oRMR0//AyKe6agzgfUxn9+SepVJr17
mp2dM7tRL6HDfRhocXGb6erwPoleFclxmyys6DgoOx/8SNno+xv0CFO8O2Kgll7ewCZi9PNgxPqM
xvuj8Eyyq22ykt3mFjAQ+eD/V/5Byzy9fZRnNusqBnATAYqxy6w4ikFoUMe8Pa4SmkNonwWnc+yg
XwKqNI+kDQnm4xQ1e82mt57Vp9+Y69BztdrCf4VLw80njzt5blSABRmPJPj4swXPtnXvejSieXFm
kLSibIzcm1xaLoKUdXxAnZdLldCwhRIGsBRLSHkdtcbfKsnQK8y4z/FPSPBWvGKOi4BecBIZNL3D
H3MpGa6w6g+EP/NCQJ9lbsbxaUkB2FEaCKe19+HTKBtir4ZUiLmJlra86ZGjPg0h/2QUnL00acRs
FZCZHWSTRVQEB5Xlv6UF/ksRppcsxMPAEwlqH/w2ElRGTLhG6gnRhJ3Ioy6ISjSZVuBL2AqGvEeh
CYoCbvZ+ZrWtcxfH0spPbhVI5Lm2CEL1NnxJESt1jBrc1uZQ0+fFNviiSkCFBC6GjgAd0kX9SQC/
TFBibsa1k6EEMbKL4zZvQSJIgqnt8/saw+UqX76E/U+78ubjLrJkxGyi+LiiS9PKtD1wf1HsdDFO
QBBzPZrzHR38kpcxhf+qKRZg0YX6hA36kftA4NyDY4+mOLT8qThsDwdDbij3bvlG9AGNrBw2Puhw
uOiS8vWHQVH2cDZuwUrBN8pwOFzOPuLYLzh0AACRuHCaE3tVsjr2pRWCpcU6JcouTMAvLPoaByvG
KP0/EpooDn4MJIhEPB9eLohlcxTg20diJ4xKYsrke8IwfZGPTdSiZrEZjW/QQbVh3if4tshnNgUY
Gs0PpZ0u1mVLtlqEya1DUEsRBG35uN+LIKYxb1dsVVvzOcc6lEYu2OEsqgXf/aAkVNraIScORSPd
WNBN2no6MqI8w81PoB4bc6HVR/9xu9LE+a3ys/gUetFBmoeX8TVgSlCfbaUSB4sfb8MojEeBqoZo
w2KXSnv3XExbUXG8v/x0T1a0YTw6fdYwQ5DLjcaHjwKFHcjHnNuEpNPvfADKT2NLzYS8dw8tQ5gD
2ncTTaJuKbgGXvUo1Ew1vxNqidqUwNfPD516H+jrsFmolb6yeDFLcqCMJvuvE4VjvDdemOwcKfxZ
Hnpdn0iTvw0Rzd5C+sPKD7ES+ABAAR6TQWlIpLC6CgCThmV3V8RpozDAy2oI3BrSCbKNv4DtLJ2z
Bz1U9teeTgOMZCco6TiTUx+ajiaCn67G0hnriAMxpXB0miSdGp7BU3XAIITsKj+Av5+SY3lq9s6W
LWXqzHHtXYggdHlaKmIcB9baOQ+l/kWyX3196AaRN9idsT1DCANFRkEk1Wj7pOTN1Ud0sPCOkvEf
YB6JTH09vLYW9O1Y+W59NTZufzian8Pm8X+yJnKIuqfQUgMxrUjVPN2JqeyMzeS564e/JkJNzq3w
DPztS5lyxEOJv0dKhbhxgmUEP8E3SRTB7asNC9+rEJn4GZSbg4xyPhflMV001V1TLLNHg30/SK7K
QKBoGp2+KMkJEju0is7S7bvANywKXTg28EvZnIaf4dgSWlrzbF1ua/kuLPBj5MK4dSIX4553NibE
9QtX5eBjiOOzEPO9n+wEN30278/ffrqQUqH23OS9RUTRLbT4fLe8KQKIJN9LgVuTtCNVg4C87pvt
iN8i3NwFr34qGGDmuOEAFqSjWNj+rzUzkiC7fDfqRy/bLX2HK0FTeQ/L0m6reyFeT25Uj3GJKXGu
vOKRzaNkNk/EeFjncQw+umo/uABVHxVew0Nq3UzuGEvFMeIC8W0ABseau7E2z/hTP3e/mS6Y31/7
rZYnBqpMEw8Q5fpWyVgeF5Y28gUGalalnURGOQBixKo79Vb+ngyBz5gjgd7w2hISPSNywKK1Owkp
8NCrq8uVwDn2WYHsMaiO508x1FBtEy9GGOKFyIMOSyksodVz7OFQZFD18dYhr9odLpYl+HYR3R+z
JOvpqmN8dDbdmBQeK/tugFT0R6qJUJs4wu0vkFL6zqqzhEdjTRk5/Bg0KDZgoz8sGcAdvlh2EPWN
9//z8OvN4fgws+yp5W9rmy57O1/iyD/FxGGDS77OoxBOHZ1vQKRbeJp5FjA0tdtHnVnINkwo6K5K
5rvbypyjXXWal665+OAFf+RW+3sJ9KRx0Nd7zuJICIq5zTX1KD57mVyuyD5/DqmgAZfIVLm4fInd
wsoBa0PBwBJIi6qmYgmQHLUPcqcmuMwER/WNoeBbGO+w+H30EAPuN2F+EOa1U7zg6albfkC+o6FH
SqvRvlPgafTpwj35vsh7fvILd7kua78SksLD/legzWvANpXmj3HIuB68pCjjdvzYjZnr6vURuGFu
49PwpauzXryf+09OKLuJ9dakIhOe2zremN5Zs3MUh2MAEqdQxJ+oEy6WAJ0/aOLZTuudqk5YL5vL
AbLFqQW0JMduNLdPOpouKiFJwAsKLz/uVt6tqXkzRhkYsX3KDw+ljk/8VULuoZtzqGL4gegZ2u+o
A949bTzDPix9rz08f5N/WRdiHYpb8nqRf7Ndq/4jKk7XMwdGNLtmMSOXCY0mkPNousRnJ1f2vmzl
WJzDwM9kLo6cZfebLGxu9NAPQgPsoluCiBtkLLvmOi4LB8gWFnj7iDRC4lj19S0VuSB3qR6Ulfr/
oFV/2JpHJ+kqyKaReD8EbPsGuJyieV1PZLOB5X8GimiyZZhy0sZjD+Xv371P5kVUvfdbrXuuiRny
o83RF/s3Z6z/ViEyCJkd8cbG3shZCBZVVBj2uVRNE3/0/kC6KwO8Jh0RQ9Sz8AA12XJzcbxZ795E
bgpeiCHwuIDxjI+btL6S9icVBndoAXcW4EMzDrWE0xkZ7WN9YqSWBMib+Im2OM0ht6aex3/1hJBF
wYVepsjebK1M5KkLfXYciRRVLTF5PWCi2Z0T2EzlRcRDKfCo1Ri7XaE+hGDFPgKhYrcOzGXRSH+p
r1VgdAzUxQaWIVZm5//yfst8hpPWiyxjLTL05tNSuo4V7j7fdDI7rSU59wQvThIxnk4AyTd7blrR
dXBEOoXxxPI/xCrqEyImqFK07mm6NwfnPCk19ILK8BOiEGsd5CCV1qlL7yPw0N7/NOaj+xYwqIUr
2pz0lJbXM+yQhuKGsmI1gG4i4+Scc0VLs4RSjp8nitjUSf/fvQSGzfMvAdzTwcKDz2Dr0djpIsw/
ikTZHzUn3Xgvx+k4xUfC7r/rW71YeXPUBZpimU+0XdWqw60PNJ15wTW8I+LsQzCnLf86qMvLQuLD
9njc665dNPZmZ6qVi6Sftg0I2R5RldSNapAkAHjRML+Y4efBVnoIjFpgwPhYzEKFdOD8/E90piHu
veeVgnhhQdYjXQqVspt//6AHxfjBhQz152/O7lSqrcVs7FJALMJUQNrHt/aJMTWG9oyB02m26b4A
JJlSm3XaNBDsfOq1NAfPuIFjKOQnrx0TvDrKuw6PQANfezZs+/fPt5aMT4TZQDKIEfeHNNlXsCRz
bT4DoF229kyjElNOh8Y3GB2yzqWQGVZQFJqAIKKc+by2puPHjoh7vHwlYt9+YvDH3q4nM9E1/Avf
zjDGMA8dLAIC33k9NVtReFUjMVUu0aL8bY56VWycKv3XzS/uHeX5vaKpBwdkXFx8VVBQ6R2jlArh
Tu4Jt9pev8wWHqss7vVjov4tlbcJoY+48w8VCS9JKNP8O52CpwyrP/c5OaJimombiub8NA9OP2xz
5X9v61GP3bEzJMNYl2FhkTVjZMIbwZ4h7tQM3avfHU5HYLaxqbc/ZrGjx5TcTQAlsE4nkDnHJkeZ
Uwj17/vW4g2o2tque94geMlnDNA6IDBVpb71qG7w4chYK1rrX0Tfq+pWWxalPoItDJF/8L4fwFa4
mx5wfsMfQxCFR5ei6N3EQ1mdNIMxMo0NHPsyaNTGA6vU1DJCviWwLtlXIZvH0w9ASBIpkcHcyjkj
6caXUJzg50NnOmdpgglb8NOeNUBNqYNm9XkI0EsJUUr3gmil6aDeNsYvlMEqXT9CrjHNLwfvIcri
WTkFz5LznyJKuNnndxjsCG/WA7ygBQrtR+lw52rzjAUt3HHN4pqH35Y4VpuVjsxu+z2wjkqSRKtE
hAWT/79mZvS22uMBQScx8fACnAFTGg+9Qy/3HJSmzTXd4np2A0PYFcaAanjVhVV66eCeSno320YO
QM/5DsFYAH1j4HN+boXRsYlGf4h3t6kPoM9SKHgHDPDqcpsh+1Xcl3t6wJHap3oOrb2YZiDEl3pD
6iCyUmgyKbCIlGajCxIUInPND4ldVaXiLDFckchJv/gIkWX2uVBkpOAhOzIZEr2LmHZSvOJHqhHa
mV9e5vaErbVSDXcVG7BOMz/mojZr5+2driQD61bukZST+tUN5mMecKzXA1y7Chpjk/o7GBrd+yRr
KK0fC4QUNMJN4OccCEQTxnt5VsmKrUi1C23TWb36xI+jZvGbKpe14YTCcM/3kXZf1zl1nNtxB/6k
ODRr4Ye1sWc3oKkLaB6+N258785tf/N1AYTVi/mlfTTquhISJDsjgCbSCXokYJxchNdCJzH5/2Qo
LQUjbm2Mf5mxDy8DVXY6zHDkeRsf4G7XBaYE0iawb3XNMmTK2sRWQle+kj0K4NrrPv7EW2OrzI8v
kt9JmkZMRMMugMcIMoGpfLgN4XrvNfyCCrVm1aTagMCkW/M23L0B06/oZ0Pw0Sxh3hbaUAM+eLym
b21AnqGgfLXhU32qYtWRwl0V0fxSt/nraxH0XFRZM5wRM8DqP9Wh2AF43sJC4niRQaB4FIbWBgbE
HGi1Fz1MuOvhIdavxXPZwsAd1tmRMfOv0EMV1oTV0yTvwwqex1OuDCrH11lXjAicoBSc7J/TAM2/
n49VtdNyEKIdQ0pzfzk/3dnkf5+Qif2AnRqxhrIg+KPASGxuqnm+kzwTsZvXmsMa3fzTX7MV/Jiw
PNkTcOw0DXM2W4JEiqyGSBkthO3KizEWPG5chnMX1X/Hx5+2a0MdrOxWdi9/jyivVl2LlnQeiX8S
y0WPcrqQ4sPKxCQCnf7bDRH8NSZuSKOKer/LpQvf4DaRSK5Ivz5BZGGhDbce4bLNC5bRlo+zwMIv
hWwfS+T+QvMvi+CLxOvk7XhumY6cNPcKuIy5HWmNwjokojQQrCKSdHl3ZOTEekgymeCITK2cC3ts
kcKURZ4vdkEPbTlKK2k3L/3d8sQPF8C1GAkooerjz+SECZrVtBQ5yX+s0EEMFJX+zxXppNJKw1iJ
R5HZ0mOpQEDag0TXab9fXIPAe7wFoDk5BPQQoD0ZWxKhsa03SmiI9gzcSaWtFlrA61+uIK5+OsVv
V8cHI3Hie7pbtKWAzEnuHp7EU4yTMRvp+uhoaTnr70V9V7Gj9SrnBA5doSwKi6Bq6YB9vv9qxkaA
l9D9uQ23QHtRE7zrf2PDDOPWWH+E4Q2hrYr3ZCBIWNFBt2TtzeXrA0qJSZL/dEMsWMhOhOAqQuAy
qb/6NBnfhA5uaONNxmRjqKpJSH31ZEzYmrMgpfjrB7y1ludWz0bk40ZJAFTbNh6Yxa67l8i+v4lS
pUIXenDWFEjFSZYK15pj6HLGcUFsTwjZ4M/CNkQ2bW0jMRW1axstJAygpO6wtL91k6QmqYuq/IY8
JrBSISEf5+cgZyhK2odupcvtJ5JsoM+MtSyXcSc4VpdB9jXpmLA6SKHf2rIt11h6ApjEXMcilMB+
q6IGtWPmnNTgLjunFEy+MerUseCyjmjQJDP1lJVOcfqXCUz4GylVuhydxGmy9vdRw7+MTmWlc7CT
2jNaAbtDpbRpVU8vKtvUaqx6WS8M4Na2pq+eLF5F/tEt4VplHJx3/IvKmIdUpzKj3lktGrG8qc9N
P3fNPt7mSDOGFP+8wGZg1V93O9iMcZyDKfPq7J5uLAgQ6hT6VIniVKUtFGjXnKjcGxs63/Pib28x
YQD1rGKCyW/wufLc3Pg+ijVjiFsPEat9EZ3H4FE15l1Od4qNXZo36A+UlJeINIccxGw2wjbO7m5f
n2ViTGoCxm4a6tT5Y0zDYEbbKyZmctxgFv4EP8lNVNGmFZgDvRrExJ6QlK8sIvbks54bv9+b64xo
KN+Yh2MTcLLriv1+ObEwd7cBhWfdbQRzYsCgDJZYjC3D7ABjKLuOiNqQZZNZHWiwNsq/NaWuvO02
6f1nl0RpSc2KIUv+akkJLJS1SS4VdXG/m7JCdsh+nOQLdlGuwv0C3oz5UK381JqapsyO9LFb00Z4
i6INR3RFyXGEeJePelLyx/4mEwzB6RVoS492lpRuW+s+PSb/seNlkVW9PSII8F+xZVX0PQ1pRn7p
5MT82bUpVuVXDuReF3rqjwJNfB1G2atYn80/jt0efGsehNYaGV08eEHQDcbG1tVfCMV4ke181Bxl
zkaNBKQeseF1fIEt58xdERNHagJYtO6CLb4yu1/pMjuPfTn+8MSp38OmxhiLfoiwVBNruefk5Mby
0m9hVyitpyU4RDOomJohGiIGLcplCrMSNlC7ved4+XQguwooltaYNAeN9eho6g1KW6roO2ZT8v6j
Y/oyDanN0C2Ztzer4scgpeLEQZfLcHOpxqmXccKfpu3KebHFA5dei/7/h0WmGUJE9R4KUdCr1geP
gM5dn+uKyVi8ao2Fd04JU22FBGvz+A6odn8CYddL8i6HdYOpN1nod4ZAjnzqOW8c2Ld50kTV/gOv
dgjjItTdg+4jfZtUrKPI2c38FHe9FKhJrg7ejceyaGTIJzIdn9fpMepxIdOc1j7aHMjOBMmV5QbZ
c21rU0GovhcqbWeynTP3I2oedQAYFvoaD9uD+RyEpvX5QUu/RvOItI9EwXBalI5YYZK0OE41TIqY
jV+A1mx+O2NXwcXr1LnnqngMa2DdAH+I2cOnxZeTQkc1INPt1ii5cIx6oNobo26sdB00i0t5DKm2
wgrfpk4+Cm6F4tjuqXhSBYnMyT5Q/X7s8Q0QmwRFVtztX6aXYrSpMVLEnqpg/quXXa/NYPtDkCpY
YOs7hvyd7sMv9KoOqAEeBFTQT6cTi0z/eb2Kq1jJ8ExLI8G/EwrpNEfHsIdc++rrcoKvbZlYhbQ5
lUB9hFMJfbBk8U/oW2AAUsY5lY45qg+dmqkjDRjaBlBKMRKs+K07HxmP5nCZcOKNpryfojRxD38q
iR1klrkg2NtZDlhTI5SEqec7VSlP6jSfyYkQeIB+KEUOrIt1TFFkrDFZ4RzFZgorBJJqma8EZGy3
nwkvTWT6ToujX+d6w4MIib8jORIHjT00HrZkwXKZNt96A8Gkr6NG1jWrwbsi+8PcMBPTEYHDa7Vt
SRJnY3qhq/k5Dw4Xc26taLJCfBqVQY7aZSw8aZObdxHCEa64kG9HjGApr1+TXU+CVuYi2mQ5QKdX
/eZ5tXT9nKKHDD1dKvyAIDDQWP3jP3yuJDFiocoxvySCSNpLI7rGP/uV74J17QlqvlcP4bXn/5Ts
/bdCg1Shq4yB9hntKCmqDYrzv709PgY46NEgS+eAvsGq54+5ruxDnRXgmna2OqXOlNLHl7w6dgSl
Ohutfh1qHOS37kSCyRAjDNFO2zg+Dyg53pZTkizE/YmKijLmyjKSneY75mi8qMqr59wvf27Du9I5
U7WKQQLg+1Gt4tW2c+dWWfCU+URwe5eZcGbc4Etxukf0jMO8mue8ift2mV9uToeOybPG9c479Ddh
eosTnjomJi7JnrrBXiENuUASlI9ImKiXM0cTnp0BcHPTlSSCDbziJf3QR7VaCCOwZiy1PBs/DhMP
MCwnD8g3HksG6SOEvtjhAIOq567FpveJYm2qqy+5zvKny5X1lvnx4D+8+swoUny6E5AKy/1KtHTm
ZPFkheWMClMWguVQEibfidT5AZAaeU0LG4CAkze43Is09hFQ2DocR8toixezb1LiuVOwJTF3vN/h
noCs7cI4AinOFzLV1qpdXtdFhjYPZEfmWKUdSMqwup6NrioJd4e/mDFyaWKhS50mLMHwQLpdNV9N
LFLCFVpTCXDhW/FkhYdAt7qCO7740tU/DlSXfZF+nmVZfILt0hLr2Di01FCkoOtjb2Fx0RAK1aQg
BkE0TJS1b+JRrLjF7b1jtNT30nlHoOKic9pVIbCfyKEcj3wsPSAgfkUr7axNiO9Y87Jow94j+rys
Pmh+apjgJFkaTYCGZOjQ0cGNxSM/X9J7pqKYQbSjBaNe+OYKUrhWtSfbJJoDIMsmk9C9lXCVLtxV
xy/ojmqFbsZVQzJSHNbPEaZGlu22zEQMzdOsnoSW0TA5OHKtQoOecRun6por/puKfRUEYBbnBTPB
b7DM97NXJ3akPHpA5smzLcm/49pY2Ju1axJ3sW1wL4S5thGWzRRUZ25dHOs7c127vXpyqLX36KLK
bfiakq+YlANwU3a+nU+vD9cnEJS8VdWrFKhc1oGqgS+d8i7UK9z1Y7eMXA/ZDIlzd/PXoYQJXaDz
fnUE+/d8kr/FH6ImLfuVlxmMnB2d5wQvukId6epsh4BAqFTJOlnViFL1ETcfp4Ik1Kgdf2hbRk16
I7Jhu7iCb+EZ9ettGuqAUPNpBzv55axV9ZjfPn6H6CzysI+Cdsmi8/plANcDvmaJ+Aw5aybaSdmD
DZs4qkoPj7jmiJJEXmxiGKyLnsFPAJi7dxLtOI+dS+ka/tgVlcUgzcTl8f/gjBd2E/BqXIOvx/jj
Q8Sr++icFa2KIYC1mC1+pEmZL2NMHEPa/yS0xTaYCgzgwn60I12GkRAfBo3vIKIJkw4C9bLIVSNd
4AwrPJW0q34Qx//JvOv8Z15HhgWL56D5ig/pv/GJfEMzolMJX1nFeXD8g1NThzqq0pTjnyS1wexG
StveCSmyGnWgT4lXt9useFN7ZW4vUiiAfpp6iT9TOrr0qzWXJI9WIvSjPQVIaw21q49r0P9G+bBn
amdD6/7xRj7iZVs4HlxBG/Bvw0jkTbg9etyXHHpYNmURiCFf7zU+9LJmFQq9y0XR93qC1Fk/b377
fXVCE+kiyXL7ViDz0MKq1//fv5/I3Kkd2y9ydx9ZEkpUQDa3KiVV9OlBC3Yj79gAnSO0lSaExos/
9wPI30eGDqlWI7/pB7RHv37bC9Hd+Y8BNuqs5Imara8ybnr5qwOCrVr9C6JbnIHzL+ZgqipMv7zL
mFALZ6Dcn9puwztUH+A9uAFNzr5prESeWYLAtVEfo/p+XZy4vqVktyQ9MTwbD1k+x+qmakxzOqfB
cqFc0y0Zd37DZwJRgFlRQG1zuWo9wTbAbeTpmCm2au02NQRsQ4mpULxDY2IIGikH4hKS/Cj5eHEy
VFjAE+q1kA4vPKHZI/kXLV1PmNskZCtGigIQrUBmwwOdxaSETaZikm3KQaKE+u7weVMhdZ0iUUvj
JANfSC7hnd4jdPQH8eMSCJXleHGYxl8QvA0efoYwXa0BcnlNzYpv9DqAs5MmDdyvDTZYKaYewuEU
R9LX+jofb80eCfj8HxBm1sy+eMBRoLv5Yr10ldtFCq6k2ivf4G97Rol0iln1wooFRfkqlmRa20rw
pqDq/PrqzPpyAOl/fncZmmDRVzndWf1y/WxSqPxCa+MsBi6VGVBX8028beIHogTOBY1KQGGIIb5P
9RgWc5JdQA5oP4sN7sE2NF8rh3zv60U/ge1gd+LonQWXUHf9mhOHvK6ZR21G7fhvVfwuqwdSZ96g
Y4YLS/PBaMtXKEOVMaqfSqF4Wbz9OKu8qzSdWZVicwTcccJdJPmMW7xzjTyGxSqH7kKrQVxz4Qgv
g5D26p//mjhN5U2Ock0MQJdYh+/T+jOWXDVmuYBPa4yddLKb08plWtagxq5qU4r2K03w4KgdpHFp
deY5nUm1aGlGiaJM+lwBYwwry+DtWHDuGb8G495nyW+Sznb4f5byb/PssNorJdQnLojzWfmu88li
OLE4ZH2TFQPE0SMq/TZFd4m69/MXtNMkosej2ccXpGhp/jfDfJkuO0HeQyda7X/vLUPa/iYE+pCM
G62lEMdsEL7AJ5/f3Y2iCxclsGKouptOcXzA+ANKt8JJMZUGL4Pyg0sJBVJxv2gRba0JxSt9vbNm
BISzXqYY1LSIYcYzx2mC3I69eiCl4eGiJAt07LEMvOH7pKzED5Gcb/N5LsaqDzuVOK4Ya15VyOMa
wvCci8nAFTHS9R2b9cZc1R8TOrx4bmqIV8I4UXSXSg/sdprzeb4wcDgzdBHP/MQ21xzQ7OquiE4T
dZq0kzLgv/ezEkaFv9AB6YeWFhGV5v8qum5fmNOXZZH1y9rzq87d/zLeku0da37zNPZ3TEPit+RM
NbtTLz6Dl55XjwTMOcdRAAupBdCjzVP9hrQoh/iK0gPU56S+J602HtORdHgAlyQ04OiXrh7VgHS3
BgV7gv7bfNR/E7ACWt34DTP2gUjUHZ7/67/E0lFfYOoeiuNqXDhInlLGqZKjhNdOcBnH1v6CelXg
xtN4VCKBZmgZzSMy0tLp/d11mrVW7Bo/SBjIDzuv2WkVVCZ/+FOZBT7U8FX/GQ97swikEyST6lf4
INKcrQjQkh4ffi+PqbQlxKQFUUjioqSeNPuYqdBJbCYWBJAZc3kn2r/KsmC7Gcbxe5QOketlZX6v
5gf4qUy9NUY03apiDWaBrjHt1bz+gicQBz0iqs7Yybn913ebYu3u10ueXmYjsUJd+uml4esn2x5/
J/wCsfGZTHxJq8mY1KRgAV/uJgU4bWs0z7nNXHrklNJ0b52GXces5uBZRd0pfu5h6xeoybVsDoXK
CkbzcwBEzm4bjPDAsUH7XftmUJpLzZ6XcESTDh29rMGCAEqur5YrzOAUhRZBtf3uIn1BeoleBZGy
AkVoeyyoLT4PMhYoC6cFDkbgLHsxCI5UjlVyOSGg/HMcT92WV9FdaUcLSz97xoJHSURJZ4S0B1Xp
EmUR4gsrhYIddCcobNGUEOGSRrMf8LmLFHDzeF/VJQindNyX5LfAYrlt/7vi682nFg3VkWmIZ5RZ
YPXsqvSZ+Pam32RD5lmY8wdhbrYvup6HLqHY2kJDacD8gdb93padXMEuA24bSB8doXud0DrfyP0B
jP8m3/5jO8zOQjDC3E53IiBJ1Q+KrgLu0JtsgS+1TxrupDUjwp9dgnzRMVh+J6GtNmbmHlAauKyG
8XjAYJU2tLRiMD1yJRC0nmek4He0PPFHVeSzkKkGuYP0Smq12BKDWdxjt+La8T0S0SlJWLhoSiw9
Xslb3sBOvLJtOV2TzzYTqsewC5UC9IjRfs/ezt7HACEaGA1dyn62AIF+WPNSRbCHlQhaZ+eTy+Z+
TQiC+Ik5KTaOdwmysI2sIHcI6NBuCT8eH3suBhXMmE3Vxku5E3A2chAi94uBbf6jYotmjUqBeK/b
wUMsQLhbCyHfM3CaRgPq2NuKHy80wxh/L6TzOXMZYjyfnctf/HRAdoSo47xWAjLod+ibZFkoIRdp
fT4DcPIitS9JH8KFWs1YUds4ueOU5q2/2TTY9n/7//KYIFAORANmnqAedD3E8HaYDE2/DPcNH5xr
iVdv43xyXwgCUYBv2zmKnjLQbTyr0o11+1ImpXfh8OiOoQzkM/XfD6iYB/UH8QPhjcS7dz5VcO11
S4izRYhmqU+a2Rdv/lG7uxmSSCJWlWGcFH50agiwSavZlLj43wOHznwKBXJn2OKXo3D/nBBnjjhz
JXA0cTSZ35GNmGQ2WuYFlWAF7Ng+8sKyk3D8/mwoTE9PR+g8xEIOS62SCy7LTvwK3ePth61HqF3y
H8A8qRAfhIr7IDuTsPesaMPabd90Vdl846RObG14BZywGwS78+TSAq7F+QkcnFlLcmodMDjywA1q
DpGAbJEg9ZhpgOyBCuPQLOa+q3vjq8lhxIM5Oc0vT1oYA1zzksgK7jcYhinQvtg2e+Jsov+FWYeY
0DGpKs8olgQbz6VvtP8D6T8q5AduLdAQV9ybaLCfozoQW0FRPWOXtfq0Kb/lEpz6H8Z3+i0BL2Kl
GYKpm1ZpthTpaQbvFkgJJYWcRnALfW+jDLtvzvaOIq7W/aPCHERfqVvuWuJEYg+qgOwVVjcXzqo5
1kuyBnq6kQ0RGY/eTNW5BVz6J9nX5Y/ao+oFxEjz2tnymo85CE+N8243HWAB0nWEwa6RXUVl5W+C
EzzHavCwrYsx/cHUGp+VH0+RnN9/fTRWBXIZz9s/y+Zpz/naJY8KKd6DZiSXElISP13/3W/+hBkK
Gsy80SXx6pBPnPVh6HW7fgPbxwJngFtBiQYjXvl4lE0OcUzD5OinRsCKb6gsNtxv75lyFT6GIDsl
gS5Xdwb+KLJ8XJh6X6A2Zbe5ow8d82IM/OOT7R6iZe7/UeqN/v0oCerY29hOVWs8A6y7g+zB5YZo
ryILe6A58WNi805OjAk6lUqBk0kPMsRLpwSzVsBuyFQ4uAeFrcAkwPuHdbbAa1rm9h7/B9h3pCxE
ZP5BoSGKPLBMH+e+lwM7VjiL0J7eck2Xb7Y/hgeH9bTZruXvUvMffmoCTOynSyUtUA7dUUN7EJ5U
Xf1g1ifXkB+d+BczdGtFcFIG6gMZvz9NULh67de9ZPrLSNPGi5NKoiPMpKi7QRXiJcxC1pk+L+Br
M0Jo9oa4jEjgP86O3an1XQlYF2VjETxGrTmmIOE/MGJuDQEpUC4K3aVRkpvCfc9HYScYjHO3E7aT
kUO62HLE6cpD2qPE6U9EGcYryXDHMibhBSXeYBBOT6lnKZRW9s4iI1AG542fWz7KfB9lzVdyXoK1
PftylI76ozgMzQdfqwarKncoOuboep0Xbehxphz8q8ZmuZjKkCr2/aWxtA35VXn+AhTZXloesSyB
YMqfVJZ6us3NxNXT0VrjW0fLn6swl+hd29PceTJIy+0b0GkNCvprbamuJldWW/ZRL+ldyyqah4Gj
q1rfk3FuSwCvs2dtJSOYEcIIZdk2lX9V9aumy7zjMLAzgoLmMLYS1lSn+wjZMosGpM7g7rma+Wtx
rpHWdr7W8abdtu1j7WsdPdH8yJkHk3zcGNX7PVJHVY1rmue00A2+q8u4KqSMalioYf3TRJZNzZ1B
ThQlrtE/S0NwGhYkp0BUyLs4vx7OwXFxcHJCIt1Nf3aS2WeAsQBSXWs5AQupYERZ0qlAE50ed4/A
JfWdKHE4cBG9YbnlJkcQcx5mbRT2o+A+R8eatv2Q3/KcEqjy7CmUQXFP4ohv2oYSE3TUbuYlRxtW
Fc9DgUutR2xRFRD/bQ4960nmWgIhfAwNtncI3XXLXF+D9lgyNcnkAgo14X5K0iS+uK/inj+0BPDs
J27jObzQNh4kdG4G1799Y1O/bFiwIBhT4Oi8WfsH//vT5uE5iQ5OCwyoLORc18sKW4dDQv0EfLbq
JhRQ4ZZ7+UJZiICkcLaF+Pv4FMI57mmtgG+Hjyy6XnHh+vPh44eUVxsQYox3BtH+lf3zaFc3lMtJ
yKfiXYBJ8hnODTez8I1+qURA032tYWml3d/XvX8HD36xt1Bf5JdF8bBwA0zbBlg4J/zs1TOxOZzP
+F3HIZ1ywGTOH+J5bhDuDSUT7aw5kthn12EpYyraxCu5hb3bGQGcPZIa44lTVutNH101XcY8Zs8J
Dr8wPXzMbqDXxfFC12KfIMmqccVrevwxpQN0yN3URRtCCpYr7hlj4SWliElLhGtJ4byUdKROX/MF
xRrB+OZv3ksgV5hyjWG8m/cmyNT2D+IuuYexn4kG0UCFDgmuDCTeS4xHe9CyySP+kD3wER7Hln+h
IOlPIoqgc/gkgZBnQG+ewta5V3rT6sjH+tcqcltnX/LOY6nopotHVTTpjfQGWwzFv6NG0K4DMrFj
BXbuSXipwGKLkcWXRVk9CqOkA4SnAlGt8d4g6W58oVCpbiuc3Mi/RWv78Lk93ZgJo8aRgGHYCVLm
AsXqwS4pxu1ubbyOdtqUP2+I4t8C+sGRb4pQyHQL2/E8+hHejkigNQWSuR71nmgHMbYJFV0LCBG7
L9/B8Bo3W3Y6I+idzPUcgH/MJ/HUbkOvbgQ7FILGgY+Dk7aZaJ+7TgIFM/pM8RjxbqssOuZb+Iqt
f5vcr52vAu40p1+0Q8h74SHLyc+OKXt0RqaQCvsDNzluM6qIWY2L2Ee4HXwYqttmKUI7R36pIfkp
OYfLIo7ZXxy0DhoPB0S4KlkHdZSIDTwG1M/x3TICVCj3WRgRrVc7gTw+W8eg5D5c4QTZC0naiB/u
/G/f5FCtBVVHi+N7frPAdJAhKDPeUIxBj6/WyZW46qOKbMMqVXlqetH6DWGPTcSzgVdjpqX0kToP
Y6KFm4k0wFr9wCUsU1ySwZLeiGilU8wqx3c1AWOD3zhAfBFmcasu1GUXgW9BKioDUB7NmWh4LVkD
I0FRlN8IZwRAS3vtFXKEZT1zA9GuYssfqoKLkpHf0A31qtTm72wykjJxHsC54nZ5waYlLkDOLDXP
HObqq7k03fQSNE89rjX5I8rVKdw/NXjsU/u+RoJdjeXTpeliNHHdC3F2m5+ohqpz82PzXBDMjiF8
FW+0GcXyDgmvyID1iYhPkLx0RrYxK1Wm+DMH3urYN3GJVUkDFIam9D+jr8ZReQtMhToBt7wsN1VI
wQsm6OEB949H52U+3VENhHTQvsAsthJGX2k95L2P7cc2c/bVbSn3PEf7uaOGQEewlIUf7n0duOBM
mE//i0vD6Kx8yl+PlJh4QLr/jqlAgHwfWnSfnE1iVpQFTFUuD4RoTfnbHyUQVJpzqL/xf3bp54Oj
fHUnsC1EXpNAJ1SnL4XUI3xxMBdFbasu9Frx+OwX5WzS3uezh+MEkQSV0l97dA6AaFH8naY9I5qI
Qy1+LFHyV1/o5yhPdeTFF2HCfn3X5potL8QsobPGNfBKX+7W5/YPFxUnMiXV1geeVn0B4wQF05yz
cZGIbzpl9lGsTgd3Ihe+KESOWLCeLdUTC5WOdeAf6Q1Gjm+vXalXqs5xlMuE1jRg7z4QcdABltn5
ros9yaCvuXn3NtahCRclKQBn8cyuPKx4ZqtEtzpERWBMlEsNV3beaFYU1S5dg0++IyUdcEBG2Z8c
hce/gKsECuw4b/zsVfqpVAUFQl1yiTEydr6geSkbFa8GgpBDzOCE4niw9hMycH58tCtG3rfM5/TY
56TUNrCLcOlTbTNT4U7kx0bE/r7XHTcuxbNRVpMUGDH+RgqMA8kLSkED+opJqfFH4L3yWAsoM9VD
LW6f3E+xhzOmVJN4TKcsprKs+h7YIajnRORdeU3ouQQPVRTClGnlS+rssqgc0jzQqDkBgZwcU7co
Y37BmVPO9H+Jm69a/GlcRhV78lBmHIstgTjBWTRng0R4CP39HZWWrK+9u3mLj438AbxG+qhy8gOv
LfTDebF9A9OVksbXNKqG/mS29mgyXh6zc1XxYPqQzfpq8JdQTs4XNTrfd7t0C3LkigFvD1A6N3qc
nCYY1v9rsZPwXqtl0NE1S60G3HQyvRYVVifBptnIbBl59H2APxWX2L1V5e+J0ffmQC0FeEjoIxam
E6XTfNbFeBXIIpne/2ECPB9aHRjaY6789ET7ds/lb2rOWaBMnXNVIvZXXIqMaU8SuOyJVxCIxgYa
ERh3oKM4/+FACI1Omalnx/dWftu+A7TC0ilQqCwmJbMzcVOHQskdW1hloMO0QDmZ34OWScCJqEYW
GrR2jkogjDwxhkhDp2+y6bGbts50AnvDdDmAfGBLpe8OH/yMaT+Q+cIzj09jlYNABmWfwqiSFrha
DCzdXemPPJ7KtdZMJQkDSb21nmdUYjywZFt7h3TUZWrxIjCvaxTk/CLsbcArrGkfJfFGeawsctS2
KghoRWXIJDB3IzjCPJk0jS3pSuZkuu+7yQCk+nWvW41hw0KZgEIkGy7JnJVMTDXyHM+d/6VmhZBZ
QwhZyZQkRJx88t8whD14kRQzEb6MOqO24+2bIWrmZdnuyrKH7VBPG0rKIXeRA5Y4mvasQO8DlGx/
aOKdMHG0gZwRC+FJU5E1Dzeo73ai9tJlFwRclF95+lkal35F0Q2h8XArzM4q/wJgDOS79dD36vcX
/KWlGY1ubtOyAejFlVPbv81rt65adPA2R2BjWiAArohTwIzODUEVWBd7hKust80mld9/1hXHGTV1
j0JiubQQ/q0mU+yrV35Bskv6ytUVnoc948h2uGS50xlVi+dAWkrN8emmr8ADy+N0tkdOPIAbuZlZ
2PvgPegFHHJHa19vPhciLSa9Xs8iVBK4oM3rpoalSgqHs1ZJMulyeYC0PkWT2KcwDwxMxTsfbmnJ
Ua/lCuahVgEgTEwEBlXxBteIA7nfsiyyI6AChf8oTWbWi5cStxMehbfqnEg9fWEBtVm74eld6GeB
DXpOjIDulxwi5+KC9tvSnazF/CVvuojWVHAWw/K5gcj7TUoynoa9xZ6PlujI7IvViJ0NamNbwwPg
GqMNxP2i5KlKss3qwZtFyRgDacfBpzBOjBGyTMkL2aVWDi4RV0G5PsaMdXCF/Ug1wOmwAoNo/hwq
ot4jYldwgHmeV9g7G5edhwYt5dNhyNPtJ2LcSVb3jWDuLSCe5kdHx2crMkqu1YfEU9NUV+hVc5tg
1yMBnkptLJDbayfwdYWelwLGMbbF5mRfVaEtaYiHVvuaf7f+tT5wC88KWKDY7Mf0o9A5hxMf4Crw
KwfWFWZrS5RaRonH6MtdUPUsE565sIxGVJbHgEb9SXYWFWwIH6pSmm809/urTVYU8pgZ9uCv0XQK
lAxAjm800EVtq2uxGHxamRJwggUBzjs4IiY5usX9fOsOdTm1Zb0OjY6Bs8FNTuKt7hWawoVlH350
Am36twuGO+xRoEeAZNduhzKlZwahAf4PWkBplFKUx4dQGD2cJs3Q6mjvdRbCWFD+pMku9BrSYn0+
e2OTEUJ5Z3TXl5cfpnUNdJ8zI8YYaxTFFmpnFa4VDezfTyWailyOrKb9lgsHXEuWZ5SbnthsgdMC
37ZQXe5wh8lacDwDY2oswMlupL2pL2SNvKzTA+9StIbbCrDaacyTNEQfbHN9QyfXNKB8sROGNXra
GIMYo0WMLDiulySTRCUL7LPpiJu3q09VYDQpb4VWU8rhU/xF4cQbxpQG88hYQ84cRHwJy6hhWIhA
59EC5c5craqhNITbPJTnd2rVXL7bGhtFDbL6QGPJU2kFocgZLkCgy6uDBYV0j3kkvldRWek9TN85
pW4LrYRCjOGkq004hecoh2gus6g914F/J+coUeIe2EhjIl8NgThvYUSBYT5u+qk9RPdWcfLY0BHP
UaXwCAhgzD9Fk7f6W5voaetUogMiFxA8qePxzmXd3H5j+274T1/wf17t+VjsqzbfQxPTyj87U5yU
zmSnaKJw16cU2hsv9hdi+DfQIQXRaLm+KU4OX9Vgn7sIm4bzrUorJ5OkmlZba/ufhKW9pCO//t7T
svhOHBzF5CK3sf8QyZVY1flxJsWJLHqmjeA9YDnYhfWrB78p5OzfjlRxuDE83jW6xhc882Kn9llH
kF3Qqm6xctQUBEC/yv3ja0yTvmmTCt7dbxSbhdZ+OcVe2i2IkWjgJhA9pSNwIuO8kaRdDbkI6+2I
rpY6z6g3x3GEj+hd7HXoy6bEmZ1U1eR9Qhmz1zvKPClRGrBPPbwMJqEEBVmbfEmuAInjFuTN/2AP
LW2Jo94DW689ZggxB0Zh9wuHeobS5s8SoqztpRpQyHikM8kbAw1XVDho9MbXNuYImTaRSegvDf/y
9U2hgjdXLMud+mYLvR4N9OpmYai5kGS+I6ig4JVA9job3OMRnIs2DFtwl20NpRNREzWjR0Zph8Du
QpQ1eOaH++I3fx/fiN5Nmm+rHO70ilOhR/KA7cdOaur2pj4LiY1waecDckDKK3T1VlWegGlwn1fF
0iGPRc2vWvbXgSi9Prb8Y/X956bnrUagyAFFGdB2J9eoGkehWTxwPFxqSN5LplEuqmY53uLNb1Oc
guVG3Lq4qmZLsJG+Vyuo6VHirYB2CptH0E3iKSGVhArRKedgKcxVDN30M+zhMAk2XA/B9guq1EMo
zUVVKvLX2sizr8HBp8y+LqsPTiE+Ea2YJAj23Arx+ABzlbyO/7YmNqRrMKASlpe4fejL+L93IY08
2dfX5pPRi9VMvfGrGUIX+FjYYwuxKnTWp8i/skjAbeuwkpN/UsXs8UY4HmEFTsFleotGRfq34+fT
VawSIX+merSECohouytLpFQ8D+fQNXY9w7SkoImMM4SO4p1J1DP9LliH4amNbD9hysOOmdFOzFuN
bYL248w5+a8TmTAcXUectZt9WChvv5IaGLYc2ejjk8a4m9jmPUn1GcF/vIUxJe+9cZjt+VIii02S
aYqVktEFeD4aI+FKT53UogEd4mrbWNlmNTNCnQP0TzVc2C+SC7PMOcwZP0DIbOtHSsV0fT7a12UF
rsrxXWKSxFR3Jv8AxLaN+3XBge9RA1M/5oPckhdSCXG44f9FxE8MC+2TnUyUstLq7i+h28I0j2sv
mdDAYHO2aT4rJZyn8/J8wX+QoMgmITWAu1js3I3wrGQk/7P5YSO6BgeXVKJw6Bx8VI9MQW0YNtQX
wVrmSDYOH0Q63rxLe3Ty+yqHGZEm8uwATvUxS4Vng4LAsvJ5rrBxPZvZj2MB98V6AZQ7RXVhjLs6
gvecShwVAlTcoT34m9+PuGJzhp61rgm14M+SW3+i2RnCYLqAbRPx2exh5LDBd5qCHbXhvJ9RC5Mt
ciL8Cv/efbn1v6p5ON0TXUKvqMQvpg6jc/9fKcTWcD92paoOEvoIAdhLdQRN3iU9zMfxudECB1vH
PdsHpGLI/AYM0lLy/e+vqB5lDpjGMY7oBH3sZ5Nua+pYRZNP3ez4dp/WKkPxZxf8Slj+84XSSbNC
zKl6LUd+1aRfpA9C5sCtlkfH6GLEDkuGbDMTRDnAXOZrUTW6bYKH3oxsd+3qU+/jTD5XjY23m7Zb
70BIjzv2bQpLJyyOtQGjM09Tr+cyBtSAkbTzMs7egkWfh/24xdOvN20tUfRwgOKFKfyvb59nVvzE
CLRcIL4+5d9pugjVm39fDKo5Oe5q+dG81sO6Yv+qQzi8ZRi3etlIOm1Or4QbO/qFiK08K+prKaxh
OhNAAK4QM3ovQFYLWwVd+H97fOEOxnPUrgnFk9YtUM5uQX0kQETVOPaE8KqGnU0n7idO/A/Tvghh
/M0PufOgCQlyiSGM+1p56q6Bnv3Pmo8T1GOY+hh1oMdpYco4BV9NivyB4uS2zBv2tCc+LU8a3xnb
2IkezrEeNXPXLEO7rkjemtWYVoHvpCq2QrRPACVcVZMrIozgK8ArtuRy1iDgcLb7fisg17742Fiq
Yj/pxezu5YHC69e/gHbI+fm5JmXlPWisQCZGihGUb95zRWkCaKmtew1kjB8B4rKrdQwxPUVheKTp
phZ2GDM25uCVctcVKIFu7yF4n6Tbn60uTfw00AnYegKlKQ/KDOXhETs2Ej0cyVcFe/qwQdwZMQO1
k/V04UgaSFBgkZoU+37eFN9cHyNLWmcRD/r2lRqq/QIh2sQMifVUwVMTb4Ak8/JAx8y2kU+Oa1Uo
dve7QoIh9gf4rcOEHzvYaRMq9PmvKwx0Eonn2E9tCaHD+UdNpXd5PXshzgc/kiF5AB07j0X6dIwD
bLo4/fNd6qxit/R21U7ABcHS5MXjqvLC0Yl7VGPWaHENnGUnAAtX9cC928XYZMLJnfiPYVenL2gc
WqRVMZzSmT5Z378PJf1StK5k8KBjI+5+1+F2ZW1KO9tbu8DIn3AHVzpoEz+Gd24mNpKbaq+1bLku
GCXJ2stmSMVa82Cwd8x/UV3h+HM9LKVAFTlTwZTUJaVFDDApkwChtl4EHkO57v28whFwotJ/TqFC
I+bgUQqai9/hdF32r+ndPjsXHtZVTv0nvV09FGikIVDDPZgaR9/Yxuk91X1xb5Xv2vod7t9IiS3v
tiq0RBKsGCkl4OLbwEhQTM4xQ5eeLfNB3AA9SbHRh4YwG6858Y93WgPSyRijoXmBdDjfxTg8vkY9
jY4fUrLSr4img/8NR03eb1BE+o9P7hJVd2jVyiw85+snFFTzD8hP3q26Kb6Ni+9e9Ujuf553PxY4
/2zuwkEVI9ss90F5hosidHcfkjR67kXryPe3FfMsdAcA9lxmzlQ8umMG3ZuXPBNeHlrszGBCv/w1
wPBazfRDPgE8BVjSRapqdboYDzUAolvRiI9bsrb6XTgw8uxhKF4nXG9a/4f3pPfiKw+xkase0K12
iC7psA2deC3YKSjwgjwmMiyEcEuAWFY+HqTCKAQ9kogoZbjNLh3CDY5J0hqzOPlB4q69xzgg0dIC
OKZzdHA8r9/s+ztY+Yv904f+rjnN1GAx3ARuytacglfINLwN8hpcexKqH1HVgCyVIrc2ZPHWc/zH
JEAvNrOHXJVgWtdnYGvLANTj4jDqmifxaqHPPAbFyPI+9dhKb2Amrld6pyugxLcE7C4e3AbQuHff
iGSQRjv3qIGNNqthiby6nLPLR2GM6AmpGMMZx6JxnaEheJBy2Ha0rBfSIOEAE3D58ZnO4O16gyiR
6jBYbd06ylQfLtY1Rpu/Xj/naIig6b9ng7r3LRcdKpEaPXpSutIhzZNuTVqoDGZvtfGhVCNspor4
vzY8KpXFms/YJqaKTPifvuvHncNBiMI/+U21LVaUmRH8xl14KQ9ZiWyWdRvwOTnJnLNYjOSrtjKK
6/Uq4X8Me43ULoGydOaqC/QJr/t/+Przzc9DLtFau3d/sXeC2X61Jbn1qV1DvJ8a2oeA2tfSZfJY
zEYggwt+RnBe60UhhpQdpQLsfymYbxrBZBSP070cj7CWMoXgno9uc24RdFixM6aw5BCVcCBzzf94
0Ymz2rY1FvrqFJE1T9+m1UEHS09I+GpHGFj0E5FOfUxMQU3GgxCePT4AtWJ6OaQ+vXYySHa4ra8d
i4F1jAbnyV6Lkapi5r3SFbmRLjqTYguhlPKE0og5OQwPBdP1rKnVarT1N43H28y5IgpOW3LKKXeq
6774P8IrCJqtb3KjpdXPgngahvbDMTxhPmW7adYoV21wNDdudykptFpm/zJbcOhaUXyDi8shjBvx
2VAWOmRBBVHWFG+ia9RZolmwv7AkrIOCWjNKYi6hJeqOCSaceSXZHL1R8jDiyCZz8Z+4G9diaE8i
IEFk8GkRiSUDLgvkorIXUnVJHx5J4mtT4h+3a0q0nzAos3zN6pwaT9uBBrknTysM2oqGft1Q3j71
kU2B81xAnY/gFDSPueGOwlgYNx1MhOUX6L0uYMnW0ZzZp+QhURBpllmqqgI9d36GMgM5L0ozDSmP
zzoXp5dnDPusuhPxLMdm3hJbt6jUpdNkZJbRYxamStF/wIsYmfxVV5BqmE6DMDddHrDGiS0hmpBm
6bepjj7suDfZKF8gG6NWti0p2J/lq0m3plKsQyubNJ/aeFiqKxnVAPmMnmvwy7SztbfeN8Aj47Cc
dGt0Yqat+0qs5nKO5FaHkaRL7TJVnZBc7VziCgdd4hDzPLv6p6cGZpAJuaiCQH3zW58amchlczu1
G9naIcLRcVWvpPFidOzcVv11XhrgRJdQfvJpZ+h/b5j6a3ErTizxziW1DezQSw/yjWjOysUChaIb
GRl/FEDFNhTvV/I1rtR50GNMY4I99fiQieU8YbQS60bxwjMkd9sGI5SHSTdxAJSY8laqGt3reI8T
xVbCt/DW31mw6xjQ0Qa28qtnE7T98RNdn2vWjCRq6Bek83yuHm4JpaAiMsL5OqRZjTcWY+RPIEh2
jt5Xei4h3BE3sCNNVkwGl95pUKQKZqCerb8w6BiLuDffrawunhRksTu/KxWYIPaWSyE90dwpcjvG
yzCjiyXSRZk8269RBRnfmBUawYvd5+BO1dbPcn93P1I+C2dEM++XgKbl64E5raBpAA9JaMqHWxia
GIyBTUC6XlYptr1RrWUHMZtgeVrVLhqE3kq3VNj7SIWwJDMA5c1xloUQIhomR9klHjxUrig9VgO2
vFFhNLC0zMqUPDCFfpXAzJWZxHAw0nBN+DvSpiuBLM0WzCAA2CZKbaKfyF3R4K7MSunPm0HNJkLA
u4GCBeZ5j9XySnI0H5C55tYpzNHIKNQ4hteeWFjtZGSvwqzPunZUoDLg5LFZgV4yhw7BuDt2iP9s
CDOn0JrIKIp/vcWBnsMYdyuQSY+jBXU339e8G9z4hPU8oUfAPFWBOFsROiXDAjkJxy4HO/5r9hUb
F3PaMMC1/YWCONDvzDEej8/Bgh6HUdn+87udkXDm87E192/nKtvpsy8kpm5A8JM9GSROm54gMVrO
XmSXRcfr/tx5qB35/634RPDBEyPcBUYOlTibb3W5FWe/d8xq5+95JsuAJ+d7FpvOV9/Ai8zuGdTF
oC3QS4NO4dsEboWxzbSSRsJJlh7oFFkhHC/CbtehCmOFeAocMu9tiWdcw9Gdqxm8u4sLLHXG3kJ9
uwbOiOvchn98+Qr0ik1Mc7pQcwDdHwqdikvUw5qAlCR9pS9kMlCgP+HqdUa7c8NIz+W4yS9bYs+v
VPiRi7eLRcOSqMU1C5oyfxz0+pfUAmMEuFy99VPxUI0oiI/Yq9WapQ+Ysnk7u1C9qw5wvmSdO2xu
s8frHIpjqJdODTn8ERvlSx5QAwLTPafydhD4s0E+Jih8cOm6hmt7xTBqo0TVZg03gHaCCH0bn8Kw
HBhQGjTuJRHE/ApqgQO6FXYmbvMjqVAjO+JVqOMqpl+1RzKgWSyqz1/SmAT/rXkLpgAqLFchxtbw
z9QhEUFekQO9HK+VDaPfQSIL1XEZg8laiKaGZllGUZQvMq2hg5Lsg1WM8W6Qav3xLAnygQvz89sg
oBWRt6YWcuQrBHthgRXGNMk+HCsR9BZ88fEI2/kthj4X0HCWLLKGa85ve9m/rCi746XRdUZ1m/9e
TX0zl8vcLkYPRJcBf9f6I4lIlrXqWF3IbZUEIkRUqurGyFYk80NMZLrCsxFxHJMZoDSu/nKqHyoz
+Gaw0XT18uNLjbToOqcli+TTQcMo7WvPlXNfVOl5h9Zrt3JvR1oqnRNDmicFLNaK95qMnnaa+cHX
AKHWChC5GQarU8AifowRTnxdNvvQUio2nCzgQkwV2EnwU5KO+N+aqLUlu3C4UrWrNYjHs/VOhXdq
/vjo98VOx2b7PFdoU2hSswUx49S5FRqJkrdta1xFgHJuDXXWpnJvhQUKuwU+JVnbjaXLLWV+988d
6545gt5FtR/fILDLAwYYCRbr9H7qg7VY5K6k9ArAXos3IU9RDJzzNJEDxErr7O05dbmoUZl3de3Y
IeqdysNGIISwlnv/m7vCE0eCQPDXTNzWMKOlYtwUJyRgqO4NlCi4ypFnvRXgDDs6Z3yFi3i3WfYv
AIWk3Viie7brKwxy+YOvr+FxhWGY1yMt44YAhzo2FJKdW8yIHZoCjqfcD/SSm1ACWdwuX0W4SWol
R4rTOH/LIcyVIY8ua+UWzIHGnEyuIZjLKQ7aXw5iQfLRcPI/7X1e+TULEdDezcewiw7KHqIZDzTE
UYUsIzEmFodMtzc9mfw6a7MgWK3dlaTzyWLCY1dxAYlL7FI4oyphLD5lPYUQ3YxquLmeO645aF9v
P2f9/o8xn91WCaOX/MOg26viwCVUwdCNeJgQADK1T0YmKkLebrvKiQOVTEboFnd8IZfREVTyQEdP
PwyRpn1p4slriw8VHGPVbGWhWuTafLx9/iFITgXWK3Gbk5Ar1f5S7dHZGkGzfXdDwiOPc0YpRuV6
5Z12458IHfC7rutqTBjV1yzLhTnZYSA5NXoO2AF6AKjSyRtN9V0hNf+isDlwsfoew4xFiek/uTFx
oa5pAvo9a8NfrPQu7F3jaU+xJC0VJMut9NOheDHRbAOO8GifNazqDqEKDgq51Z28ZjCiNjy/B09Y
aG0dWEe0+HYDMlMQ6lVO7w4JsGJmk3dWH1cJTLx4KmBF2LIV950T0ijnmX7IiEWWRUqfTzisYZFy
MSIn3kVD02ezS9+ibDGeKwPc7dMvqrCcCiyszs2e97MCg1c3AtQHlsxPG3W9rp00csotrVkdoyS0
my7FHATe4JK3htzyfMpfbl+hq1Zi7xQShYNMfjat5W4wcmA9cbly92Ghi8yknwMTNazOD/aMOghZ
JS1BEgfbPA69B8SsvJ0mcyNGvisyAoKo5YWujaXcXxtnSdX02lelcRMxVsQbxjsTlnfdM5hVA1vG
QQ4Vgb0EjUclc+eVNlC53f9XAx2O6DOpylMdwRga2Oyp7VcKT5jdv0nNrf2y46nMBtTaJTPhRWRL
utw0M65KWSS7wXZq9igbG9QlyBi8k8KJeN0E8SHE1EeO6gmuLdOP7+cIfvUyRBmESGxk1j5QHIjp
BoUwyAiex9CAM0aV9NIqlrkHV/+8z8hKIQH3zTRFqjEaPshI7pEZlwCJ873Yb8sGJhZ6TMrFfxDS
0YM+3QA2MzktS6TDa2ZWRC7CCRvXzB7nxbSV8+qLSQzT9cgIZ9ezc6BbMGcD4lS/aSQEQDSa4qHF
jKOvr3HbZzvrmtGw/JRGSK5U6hb2GX8sZJygy1zYQPX89xJXRKrPscTTnP539KDuUEbchf3QI3FI
uvD6MpzTTZsOmze+Rqm69/B5cVKMMESYfF/NlXJURRtzgKbeL6v8YSZCJzSb7SrI/vpredllh1ZW
XhVfhxpKJRcbeLTzAFgG3aQV/5KO/kiQ6N+67USyMmtSClNSANZYQudWeBFK7WauSX+9Gz7GI8EZ
8cyuoXcAYwbFWVFaV0k0Sjbyd/3W1WZ+ORIT+0IDzLjv2w6I+yl7D6GjxYO2WIV01oCJpaoiCWm/
pn2aYyq/HrbzkdVtBYrP+ijaaY3PysTX6U6O8KoqDeSbA6iLdnpN27+lVkH6ZsoXI/n6CiKmQz3g
ni4dCVJw6nrIy6/hQDU01pqx7fxl4IY5QwEdxBb3cKCKYW6lu9wOy4W3NqBFcuV/1nBm5P0N0a2o
r6Lens1FaeFLeOKfCTM+rhSQHvO+YFd3kvYx/G6fjmcAd40cXLKiqVClJ86PfalY4z7bxOSv6Ve1
1MIuvsAWJPQlUlDgEKer0kUCRNjbH1DJGJmPFATa2ws5pSEh5CpuQt6CxX+EJjANFdUNJy4bQYHW
y/0W0R9CTSijn2W3fM57pTK13JB06trRNv7G9e0BjL0BDxKnw3N7qa9bf0SHy8+Wedj2AatlHW0a
RvqhDjViPkTXjwciUIWqnPXDjLwZjlpjDeZ2aKqBJLndUMqoYGmJ+O+A2PJV/8yjoA/+7az0f5rN
k/3G/xUv7QsIp4cNnm/LHqeu9UfsJY4zilnYrx0EZ9nkDFNgnYhiOavf8AwzeQN5qV04Qt07FFlT
Lryq6WUr/1gLbMZr8YMxiXR0nEB8k174WD4y4rnlAMNXFq0Lmzm9iNSII7JmmwKh3m5tMzJ1GHIq
PkUg9kUvwweDsXYVhNq0K1q3A2BuTNezQM0L+G13Ymc1C0UsJ1vuwm5O/6qBGp0sdIp6Hho3t3UP
S4T7xJDn6prv+IX13V2whf9guzkONAtiLVeVwWbqoliUEWvzIsVK7kEJIpPZaRQcjNWyKmsxbJ/S
qaTnsXT3EywL2fbQg2zRCYaoiVILpjhm852CDnxTi8HBddQ8dtH24EbY7IyGtlqKGs98PxdkhCBP
w4xD9SvJkLDZuASKMYSYKYS/PHqDQRGWBNRDN622iVJoZT6N9YzSyFsl6I9UZeF+VxO6cbVZro+Q
lxpbeMYUTp9n1olDZFPjHxab5u8KAfSoHsIs2JVw7YbJB7pE+jdWAbyaDER1zgdECSCCQFXMFK06
ARcKzusfe93YxbRJiAeAxtZDnE2omp3h4PUqCKQNn+WOSyntnQMf6fLFKjtjUHSLd9QdduWtTpy5
P13JmiiE6z+vrXM7JvHT4BlcOCrEqy7x6c+Y9utmyiVeBiDI1TL3UjewP6LXxFq96AUOIk5KRBNO
vuxxGon9FBHJw6cMd22x12tJfxE+1aIL3C2YfFKKpNjAwoQDjC+t5VsDtEIhFLdjjVFpBvSFr9gt
QS4zZBey/+PYREafj70w1lIzC3kvkwFCYeiQ6jrLFlhSFivFs1N/ODsQgYVvkYmU8o5v94kbOoLY
rZHMjEJFNADX3YcJ+aEAH4y4eWvqOjQ1jWbYhgz07oI+1E6lkoq+YN5agelkEjUEfmuCenDy5x2O
zwQ3FR0Y+AtZneETvVO2SVmuoFNuKVgVPFWVl9+HQUcGW6XYvCqUgTgDBpiJITxk/oicjMasYDYz
02L2hCEm+Vmh4HjVC4yPT6PQ0qWYMyjwL7JjKQhhYdPFG8R2oZXxnvN41MKeK+sZKCr2tnnYeMwr
is554XjVss+J3rfdw+28u2nuRjlEJyNmFnu9Yd5+gzY1wq1rZTR2RsI0NzRAtSukhoitOwWqXUR2
xbPGWdqJI0rfgZ1e/yCcZSllaPLI0i4t0acgEFvI4ggmnCXOCDMSXkuhgKpnZZgKtbOqPkyPCG1n
UBuTIMC87Lfq1+hCwVawQ0JxzmHNX5bpL3I85Jb4Fc49Iw8kNdmu+GrEIw+1uP1M9ksx5FzenJFY
zM0t1RRY6+ZBu0xbjHgim6qKCIegadt+V9RS6CZL3KSB2mrEbDZAYb8UTpYfarU1ZUV8j6TQ8IK9
7x0jfkegiilOuW69FZ4284b6SSfMJH/ocAlIffhCIkBfmXhiqjSi+8V/xRbPClp4w0jknfiQfy/w
O8m4MGFAOV0ilANoZqkNHswygk85SD4jYcyzP3Q9Yyy+kYRhd5cszsWdIHQwQaolyV/HwXRuvwPS
cd3y5w+yS+qQfsSsCxJivAmhxMKwJi28+Y7IlVH2BUF4Dyyn2eXFdyqEp5D/ps8wOoTPeZOxhi6w
Z2F0UVCj/PJHJdBA+qf5030w2Dhs5VcMme3fdBEmrisGrbFo8aMF216npv9sNl2ozBG335ApnlVd
EEPrOzTkvuwQBdgLYTVosJ00uy/R/AJhplUkqetzw2NxvOUn6/GzPMAJ/5zsN4tHCHgUxnln3Mic
w6NMyXknuAM75sdbGKlcphWfdFCkvZ6pmJRDDv7t9tZtgaRP1jceiE4oJsPyEp1FVpKO7W0Wmvck
NIovcdpnYcaC5YGLJGoNxu7dKznDBTPvJJAhp0qITwrI9JEaMJWRabJ9zw//+CSYfhd+0DW1dMn4
+k4rxG7TZGPsaUXr/DFC+66pCbYzmDiaeDqAQ2jP0eQSUc6NiVJJeuD0LEQXOAccR5udRLT6AO2y
Mr/0EGDkt8aJAm8lSzoe10w2rOK5Gcm9UnhfyfUBurtJAWwJFBP74OL85OUhqWCRvhM9JzrLsXLS
r+kI5UiXhNl9zZzGcK+c6C4OGzBcGkirtyPpqElf8zmr4kieYuCdLhVUCgDgK5+PywQSvPUcK/q/
785KnS4JxMujbgU26LRZqhRzmFrLro+EmRm8FfdiI+iAT9m6vUBAXvJuEWE3AGd9zkvNoq7tkjoZ
cqmiOU2Ju2Bgn1m6psX2HvQOO7metBSHUFvwDmMrXixfyHznEbpoSqa2o8VxQsl8xzPZ0CHTTBxW
2fTPlaFmrzXvOfzvCzVvGcqnygDUepqsBMiNKJlT2Pce2TIuOPvmueH1fglVZwJA1l6G4NG0hxPV
Kxl3HrqHzcZTLC0vb7Rbv3suulG8QN9fMBgD9Wrs0uirs+dphMFiCSXPQZolmrHBQJF3Ix8ezYIC
ODzNyqPSRHhehKxNZAYwpzLts8kXBHWPibsTCgfwCHsG5y8ghipau8qoRd5hSWoLd7c2f7/DhWo+
jIOHwohkFTKsfdumm/WCRCUa3L0u2jTP7SxBuH6j5ATsCrdGNRGGR271nIgNZXKsSFraitrgAWxK
c5p/GoU69LhaycV+HNJNO00uUxU7Z0P6T1eakoN6hFE1CseFx8crBrCo7wWXLUafxXr4cNSv44Q0
/wCVKGZKE6mGw6Ka8HgulktAqHXPMcrtInyIrJXmgcwopGvJwh6JcNvx885lOCSQzUV6JxeAKeRx
5CJ4BU+cFdEZq+NoQ9sAkUP+PJz0LatPe7vOAAiWkf26nWG21UVKqWeteCVwGmaAF4wP/4asRc+e
VKSXsUNpOre7SGRT0PyyzLRxkZN3cZ+5lpFaODw9sOFNQMAHPoYse+TTjO49TJAQrgo3EgMJ8eer
NYsSHz52lAFQySdtEMewRMnBbJsj+3Y/DRf4hWxNsdXcavTiV4PzUOPZGMQdXWGp9dTPvSCLakXw
YCMmHAzp3hYllO77p+R3Crf2FAy81X+fn7FSC324d/5RA7mtJag4Z3M6Al+cRKZfGUgMNW1/asWP
HWla93K0y+spmbKbyLuSInkhNIlL/aC+4dRvaEJ2Rf8SSbyg4N6ZfGrcbRmBhmHtR2NLkz8S3SSw
+CCwPrL+fJD3qEqTvPo2dNBvUfM7zBr2FMUVg3mEVMs6jfiYR2yP4Rspbv82fd1Mfv8QZ6nQKG9D
CFJhGkvlTT8sV4s6g9EhbhDt+IaVneb45LSpXLZbL7hjCUoq4sUx/VYZtWxGTgtUfsYhD8I9lzjw
evUIza63kXMYnJje+8cExxINgZ2LorJFjNVrpqkGFTkMTP11DKIl5NTjYtpFRoMzW9des2VrqwKs
FlL8TeyqF5xwXlSbgHmFcktmH6n0grmmnIdD1sf8qtM08tgZ1U5Q/TR4+KNi3cHu1GfxqaBCRtEx
yuoZ8PmH+xR5w5uR9itoP1/TW4kWJ5TnESnEUYF8CMUrcmxBev0GfctC6Yjk6e+lO6ALLCmj0bk7
LnlvhlLa0oQxLQPAK8xcFg29CXP1GUqoZuBBOIapqutYF134Q/0BVDdS8qZY4JdygY7Vjriy56N3
E/XVKM7WI/Yi60up8Wj9LSVtWYnnsSjjgvvKIJvxOut1NaKkqPuLffmE5mJqhfEQRTM4Nylg6l/g
yaQXNQLrbIhUSWdYjGlA0lUPznZeG/dFvCDms6cWBekrw0/gIwSEpgdD5S1xCk2RUpv+oI4kHqth
TKyUaIDUoC4F+BjjEPNhnzCY+QBP4NifSgGZQAQPeJwvXVkrOgdo8r597w3WlHEqTzuZceWFwnmF
f2lMJJu9R7sMeDVG2rCRek692HmCWEqj7nmKjE1bjQ+EkC2E86nzpJluU/Jh04y3Q83WTBE0Cg19
n5jqZXDqHy+DzZt6LybItcYTZ8op4kyh2MfCtjpUlvaMcRmkdaGs4SFCDnjMOw70z0dSF6/phU2Q
6FcxPlQ/rwj2tWOlTjNqAbt1ZHH6xJVFopiEO/d5fA0sme9/jK5GNJ20iv8HVe5Y2RMla9vBLWPa
GSFihIrDjuLgwLgi/n7yycfiZVfVaXDcdnqEVUyJjefLvEb8fn6Knc3UP3ygZuGFQ6r7kAxXCKzU
6idOsxFXXrqeLb/dZbQAaHQgL5Dspa16bPZq/RrBkP5cH0f3kma4xb54JYCFbYfr/jYcLoZp4g3F
RiVURYUJbqZ35/1CrwXBsomA/4OGq+/8Lar9AmWyvTTketatNpAcgVhLTSeLXYI1Deen0Uho/LPT
S7810m/yGb60/YATlAusDDxgM4iLZ9Nad/DDZpkNU0ImsYZICeEnXYw6jpKAfWeNE711mqXH8iry
Og8cmOe1Yr26wHBODwx7jM2/I6hMHlGaWH4ZC2B7+AEsidJ54/f//lJraLFN3VSrCCGnMV5ZsbUM
VfRzFoT/ohQUk3pBiXmZ4MjNq9lIpOlz0RCWUJimWIbEwcgJgZUC3cmLjgkzFCDz3kvwMgYfM7Qi
XZveDXs5MX0upx9fI1LCmlvNt+tuNVabvf4PadghdV7cQa6CvpHmvAiD57b3a6aDGBxvs6CugUo2
K+R/4LXy/QZMQLryqby+OlKSjb+vFRt8qs3v10b/JZJCIXe9oEzJOML9n9MoWpVHuYeK/2r5qqT7
5Id9fK1Ney6cZZqXxJrMfcfMRfQjMVeDcQWtfnG81ayEnw+Fw2cLjunSb09d6k2eajfiypVwrULq
cjs4Mwc5Gu+bJ09IJvCskVFeAgi5z7y6H5bC1uIUOidqI+Fuq9y0oCyvUDaWCjNLezSye8shJMKk
d+BB9L/L84FYc0iDixqQRkURBOXmx2v+/2iVXNnsdvhGOG5wToQSgGXfOg7cp2eeybTf1T2hvE14
hEI/wZPBrjoRSV9hd7ZWe9PEFq6r/REKDK5tEjzWwieu4VsILbcifIjZKZUu9Jnfy2aTXZEOMlcs
dRUOkYU2pi1fr+e44owd6MtFjRmpdDoehop+nob/eDXojU7EUdABIsBvpFYwu3WOnDeDIK4Bwstr
ngmIQo8UPe5AliagpWgLLnVWmS/p9Ndut5owV8NRaYDbHNnDE732SyIqRdCCh8zPhU0CpD0bKsHu
evd9Ed1L5ugRVumOo/ds8eNqPcj7NFP6le5ZcJZr84brbWeJZ+io+8qhAWfGVqLtv/7T2Jd34u/w
fD/FBxB/fGy1qy0/0tHj4E9L72CtD9kGqhg1mUEMuM5yB22nv7ohWarcoh2ISw99vtHPujSgwtwI
gw2B+3s1ummDQ2Q+bYBTVmW5pkfpLX0Dv8YyGr7hl5hkV3S02QE8/HHLZDZoXikbmY8ZUzKtN+mG
z38oEKYs9RMXqhgfzlPEvNtpiU71Wo9R82MgMkp13jnoF57bs7FO470Q7fi9oKsW7cnSwFi5W0gy
RRygDuODFBabp91r9FHVV4JSizH+Sgl0yJAk4v1dg+1v16w6A7apN3xXAD6FAmTn3pXwEZyyP/JZ
z5hMCzpQ6lq9uw2BuL9zFjuLKs/Fy50DMqT85NwnZlZdIbIHcy1AGwPwXRQ4PYIauGXGm//dyLvL
4xEiTVHvMX5s5H1k1EMwgAfMWSOmp/g6XzRLkOoE6fg3+4wAXNkTV6xJXnVSpEiyKqscmnHYCnje
ssP3ofIKr1EP4e1EjWrJovQ1AG7DnfKl/WcTnlT+IZVyvqLrKCQyYkvL5rXVdV6x0Vb1VMsVgSPY
waGq8hSplHnlAiIXUFPltQJCJz66VUjPnf+O4kMTyEXnXmWH6GxFx48GVtfd+7R5cQ5HM5JxDoCN
CDW/UmxbL5OdW+IqY02u8RP/vfIKSi4BpgWT7jXVJqBEfRbFK6UHfCG+tfKQIEKNLOUv8DA0my4K
TTdW7cfjjax3BfSQydqIuNJlY9rDKcppfx/qjqr5/2wSagFwdgzPYsL+Nc38olqkahjRq2V3A6BQ
9X18w1c2wYLvj8qktRnsZd6pI2ouacv1BFPrJaPvX7xQiDhmWvL700VYoDWnzLCm1Kl1FdkTlsuF
Ws0DNwrUSUp5TnLCwXnaP5lPmE53AepSNJ1wWZKRRuZOfXK/oiz7ZekiLIksf4I2G+MgjkTb3DAL
D8mwXETjCNs2PbIhFEj9wpRx1cKhwNxXEOkOJJNESFbuowa/GjGHF7Bv0oTSMKFVUJHE2eAHEkOp
rZHwTCPRxlJoJUcps31pO0dh5rmGjXoevsCUujznQ78N+7dEa0Dc0m1RHPx55P7tPgZpq4fN9wH7
zXIk5Z/EY8z3V63iqzdOiu4FQpAGP/Fyr6ceG/86htGTWcg6oh2jJ8omDNsgfiF3wqc0lK9Ykzn3
mlOxNJ6dIaPVF1JA67Px80atKRT0dGE0dsLK5EFyXrqsQYYUCM3qAMquicfki0ivomR/wXwI5I8a
t/Zs3mkrEtv5gfmS5CLBw5/c5jxjnSXu+fcz55SlZWrruDEE4Prd31BkRP55Bss9W0jhW2H6kS3A
TeDK3wJRNfdB0xa/S2XAbP/aI+Vcdl4KoEwpTKe2LznpTl4W0K7dHuzZ+6T5jCmYRd4jcXvAsMGM
shHyOdNT8q3fEiOIwj3ACjzwGOC9dPU8zdGvMvu4vMsMnwxGkuZgl+m3aZF2X+T/B+SJvrq7QPrA
9XMxui3p1H6OvrrJlnmE8YGDljXau5H6GT1XSyqMlC/6HI0VeHIZ+JBi74S/mYb0m+AWt0KRzAC2
1+iXNAQuX6c9KioXZRvAVC0kM7mf/YHRwq4W4fkqywIiXZ/xJ7tOjjOJWnBFG5v7D7Ow/+sF/AXA
pEkECZferljkN8qCb45pkuHBGD1E81xg2/RibCdeKyH1aVovA8XCN0sfJCO/XwwOvVzDzEdBF5Pz
5PJoGgmhj+/ILHRvpweT2EBVD7a7R60p8f+GdshWNQo5nKBLhRPGOoBXZurUSaKQTyLG0+MMbCaG
+y4OOTuyZfIVOSRWi+WDpaJjsKnH+Ajii0GMJdu3E+93px2hnv/fqVpFynwPEuCh6v6doA6dMaBa
48Ys+MD51yev/cG+4f/e06/kUmklmb3+mvPEZcgDL+ZSMeIStHqzsRFUhe0vhA73N2JUfMwpYory
uBJTA0+dK4EQQNE3p5ZNGiN8l5RRwAtc3wop6MvSlCzmrgBrIe1Gladbjm4p8fFv46Mcla66h9Oo
2f8e46JZt+mhn0yYoYSVrRhv9zc+keIucRhCxIX9Sg9UQi14cZZhqJ1mNYTm+C1p6NHpCrgSzYCP
Ng5iBY+Wpbpr0CyjUrFBtgr7xvW1SgITvWVAdQihQFpH+/5vbB/4P0Yo2w/0hsjHmOXw5oCU3Ghr
14FeOGgoLZOY1twYJ6UT6ODCfPSSJPUA/sF1TaP7+pQHGFREWN9HufiBXwv2yLtGCHUmB+rXqxMP
UMklk+NSWaVyIQeW5GFQA3B7ApElJ51MqVAAx2byVG27F4TaFHf8ecSYke+AZcqrn61Dq4BHbnTq
SzHbIcsf8aEldRuYyEsFFtuqincNXp2TI6RVDQ0PfbXl3YxQ76+5EUjAiVC2Md23VM4by0pNpVft
HWx8jBgsA8V/pi0Gtn8WSDCEKKunjZ7xYsaomhb3dIWVNcE1+YRjGQFcwdFOOrVHNPunL6wHZV7d
6swx/Jpow74+boPaWI5ONaPqLJPwIK/Mvzq6FqjzDLD/wEQmX1+WIr80qc/0Qdm4HuODOWURGm7P
wYHpBCA+EnmHFKLvB6kpeKOc4DJ6UFPXVTE1WfLZdMpNSfVeFhwGQ5ychaEzAI+ALY88/F0OAjf6
QjJgLUgHANf5qiMg3BCOeTgwV3DgDVpCb5Ws67iEKWw6UrIwfsKiHuIVtn52yIHyEXbNF5UWA3ml
TdffLa3KNvSaVz7RQO92NvU3pho5SnUADjY9FvSPpKJO4sLQBHOCz3neG3RaUA/dV4aiYll6+Y5D
8uDQ1ssufR2Ye8DpXKu/vKmTaAmnlMWribf4fU+5op2ztAevfsUDD3vkmyeuZY35c4RvpPkE5jPD
DpxhNjuDpLbw5qzzivW6LuDA1Fk2fiRloX0p3X1M2dgRQecnmOVYg4ZsztIWe4zhkzdJoXGDEUdi
vfvZOb2/GBN5XriXQy8+s8HrswtNSrLwfmpUZQqdLb424+MJGNSApy/hRIAUUyMf9jFrSkn5Q6Cz
2ckquj8DcaS7QM4xJXq5ympTmXoUF88ZOAplcy8s6OOmnvF0wfDzfACoB974SpioE8duV+D+k9N1
cn/Ds129sh+HIM3xxIW62mhXRwi3U0XmO9hJWD46WG/y30aZqrz/NjYLhC8hKRovGQqOhSnu6QOL
b497/Ujq73D6eaW3cXzRQ9wQGVUFh86tAJC1JMPPWE/Kon+UlAiQfAE0mGVFwZhrHBu46O669ZNx
mRTPGThc7KUVTg9ZL7UmRG5BJIFj3SrNbjPqJeeG+E9BvZGR7Ef2H/jHNXFcxM5ur/KUYSOJS3+K
0CJsPmgLyQtEA1wj8dKMLYJsm3hrRg2xSfKkCK2RlvL+69wW+SHsM1XLmGmSj8sHMlIrNGOxWYJu
t4nGg3/yJDsWKAm2n0lJ6W7U+RsvjKQFmmjmimepklUUUWqlxEtJzcKiW5H0yOGTHo/XEqOvvEqK
pKa+EA9aqqrOlk6+G8IG9hYqyoOAa+3qqmu5qdEK6ixAtFSAixfTzhYuK7iJG4EK7C7TdaWOHzhd
buj/A7fzxlGHlBPFmo+76hWybgXoxPZGv0Cj92gAiSy2B8sIAt3H2OyMEw7FP/L5T4++ZTCF+tdN
oG2IC0tk3IeKVJVUECihAy3EKtjZnyauvTAMARI1MM+8j+Dc1kjSLnCD02DbeRVKZu2FHVcCKxre
dUVxO8m4Q5TI1X2CtTKvhQEnIB8FluRopI4nBFe+5nNEumvN+6HxZP7ODIQXt9n3gEhe7126miae
Cbz+lI8LPgiXa2g/UUCzObXyust1AjKZof/tNH6xtGCLbkytlYWj24mCt08aXW03SM6qD3VKFwI+
vJMqG9sU7g+7vsMDMuLI6XP7PuW45mbpx42ncPdX0yZOgXT5wdwN4BMYkcYC5o8r9cwo95HvJd/+
UULT4VBswhcvvKPyndhwmFs2haRSAd49GTeZpyjHi+szda73bKdeZe3s4Kc/VhlKOuUzrWgtyWXD
naeTGUe3GHpA2Jei3h3Qca7VXKWvummsiKEnw9TYiQBRx4NIHRZ3VdFxZP2gMHVEhwzt1DzKG49r
J3bjq5dxW0uhBsIcwRIaW8JV4TurJymmrcfEbnqjjAMomWf+VnpE6Ey7AdvE/HkFlCrRYLrGTvuc
Tk1LzS0K70cVosrdPKoqmYXiiHfji/Stozq4NQXZDbqpdWXY0GCZaFvgdyFSOFlBqY8nefKq1Dsw
UV+E1i4hJaDy5osqGl1hLIuTt6AAA6RdauY2EP4SG2iKRFznsyzaAsdSfQxOb8lCsQkPWrx+rex9
+2RPVvt2Qz/SVs4lxZLZdYZ+b3olup/Vlrk+6rC6Nd5faT0/ZWVIuljws0fJZd/nzyqFij11+6QC
5Hjshit9gEKrox80e7P8WTeXBMoYVrALCYxamzWL3upg6h9nlCe1SpLhlGs0yVwdCiITZUBFTB2b
MnEW/0WHaMrdpBbWi6KawNj8x11EsxAi3d4tyKi1QH53jBT1KCIPijJRVCQHZ7MKmRATu/vRa+n7
BjWEd0EozyZ2WLqoAk5lT5chrndfNM008IKAWCRxXLXZIdHXNffL8bO2lj6YsyC5CJyDFyIFJc6c
/DupYfi0CDLnWSjvFA1DU/OWsSO0VY96oyn61WwmuBX0NFgfvi7RVmS7AcWLZ/po53YPD+PW/IPq
J9VxlTB6qr1aX8f0lhlHAGYiX6FguRf0hwJ3NbJ6PIa1VK/UdyakUjPx+cVLx+DkxJCvCk6wf9of
6l0GuXNF+DxlnUqnsKf86hxKWW1cPU9Ov9uc1RbmFs2yLuguOFXpk1IautPwlJEChDGX2m38kWPo
tqI2riSa39GjaEp5Oph7MEMGORKc6ebfpm2jlP2FrOlzjFaNad+WRfjBCNwzMT7nSS4tquGx9Bj7
wPj6tXaDd5oSDTaAkQDBdjdFSPJmHEjBAHQdDw2K3EL6QYXK2cIEGN/7XO4IyWAZ+oysJ/cHFiq9
K66VGIF3Lupcr2Ii28pwnFqOJFLBhrUBEP3pha1RBgf7hS37CFQyyh5cZvP7258HKALxzHQw/kaS
oB3bzZQzf0K3/CkWHSMLyxzX6U1HnIditdUlFhSVbFl8pwyK46U7AH4IaK1a2Y0yKM7rWu4jtIs4
oOeKuzzZQne8sFA2rn2XzpIqeuDosLWMG2YKSD3v44SZGwiSeewbRMGpcl8nNyH7YIoeLggJRSu/
ITS/z9vcQWclDbgTCLOk0KxZIGffs6sKwc5Jvp/8Kp4JlXUxY1Z1mzilgLp2p7/eRlTjigUuoP/n
18ZdS1v+YhwjD8XSVA2AoUfMyHoGskChpP3SJi7U/BWtJ25ANY7xcau2dApRalILkPtvPMuATTa5
zxbRHksxL1R97bDirtJiCVOpLux26ZFK0tbfDpNSqdhdvLalp8fCPwwBOcZi8jl+A2zy280znspm
/BJYAIPIxZFi9vv4qLALdb2ytObv5GFA7zYvALeSw7jDj7YqHU8oafani8BuzplC/mGsYTojamnq
FJ5LL2Xs81wbZySTxYTGiovK3P1GPxQsNNgLAsi+ZDB2mhy4I6YgEJnQCEv0ZSr8fAN7G2VrMOR1
hk/ju1jBK6oTabPtUlzCgC3ITBwx5/Ws27Q4MN/MRh5SXZuC38KnKjK70WThOgn1kqhxqzs5Gzye
n8ojh+tAxkJyXrDTQnXkiLxZsRyW91K1RawV8vgM4ARKCGeQx0sqFs60P7Y44yda7sZqYqgPtDuB
cyc+DUgzVs6IFMzIEwovUiUjeqjp/mlVSLykGrJ9TcULCEuyHldrHSI2jOTvcizzGm3WgOnLDtao
5+d0a/NT9OUb/6X7iBOwRpT/6ApCNzF0RwjeiXshqWDItl6PuH1R8xrEaBy3zQPs20ovLkbGjnkr
OwSBt3pz8qLHs66LcdH00a7rgI6fy/incJ31HB8RPp647BtfgIi7ApjXx7GuAkY4obkV/P/Y3e0W
2LGpDqJfnclbMoGSedsP13/N07OALpaxH/7pgtpJhoGqSy13lBILP/YS3W8KYGxO/30/XcMGn09h
V65zTzm7eMq1eHZH3vmjbHk3vlY8xku8wDQaKMbaqPo3qDFWs7l22yYW7Jg1C5Ykd2gu4cNXe6ZZ
775uf8ARM1Uc1yiVQ6ojc6EnnqZOV+jsPGd1a6Q2OrN49X7ofH/S5Fd5A+gCmCiCfW0nRWZ/RHwE
ChbKljoiV2AiDH8cNQrdY0GyJX5AjO1K3YFTodVfAflYFHYYQFYy2bslLkxIBZwxL8pEd0cvg+Ly
beQQbg4VzW56HxbN34JLfY7Jr8agXtvwhrwU2FJ7mTAMtfuVcIBd0+vHFuRd7Yr2hZOLF9YrCUos
uSltCFC04q9LtPEkyofH4qJfwKtMSSl/Nbbe64LA/5RGa5QvL7UtHk1jpxYmNKaMAHIWkKQ1Yq8W
ps8zqwyrcCjvGv9OnCuyyvDPCAKVHdf4D0ZcAKEb8SjMFt6jpXpRL+bdmPyVTb1kkCscORAO26cq
YctKCNA3VkrHFf7vJZsSHDHLcobX3aIIe/R7FLwQXOrmmCkCJq3yUiZUALSD07mXP7nMPQqlGGQV
9h7ikT44D6fxvSuHBjHX7ykB3WRsL108Y4cUIeRouv6X/K5RsVgCfIbHbIa4kGtgTyB2Vpb+NTWB
XO9YCOrU0wlDQr+q0YKZ9m+PhFnpXW98qMFR2tke36XwRulIcIOR1nMAbScAdAU9ybMF4Qp0i1iP
ScKEJxoyjUWfCQybUYH+iUWh5IK9C9YUiz8CIV07LiI18MH4BoMeib0JUtWmwBB5nHz92vj2dZck
5VczbZzJ6y8ezQ7Ro4DGCJG/AisbEcQg6E1i9YaLqktnNzs0dMwcIoTMuXq/moWDOebeGfTH3UWU
RxuXYY80tXPHjCBqdk6xQtbSW3l/87brRfUdAxdoKXhMTB+0Mzb66eCSTPp6H5Ix2gmErithlUvo
AyxivCPyExKSUu1q4qE8IFKSm4AgvHF58KSeXY+Oa0sjf8w8oEiagZnigE6JpGKSeKHQzhsiwfy5
ka4raEo8oiTzX7zqfVIMTbXNkhVt4+VMcKLxO1GapOjXADLXj7qCzve+uzCMUwilOM5/pvnZ6oyA
DHqNL88D41OcPZX1Mi7sUWpHvAnFdSSqBWcylz4ABiQGOS8bhralbzUYl48C2F2fSMlBtjkB72JJ
PZf8JGSW7hgNdckPhSq/kc4NRnsce25buQFVLOZblAQRXKlfHDTSENncWj4nCSyrgi7tfsa3vHs5
Cg3f1krA3UnOg4qnw7RTpbKiUJVs4edlrxXT5f2mCd2ajRUYUFqdvuSfKqaLYTIX7DDA5wjPaPn6
/EnLtCKYH23PgnDPg5/it7KjS2ewEoY7cjjkEpfmyu0cTL5m1AIKaxG3TYac0gKz2KzjhiBm4s3R
snM8HwrrDWod+sGpRtYdcx8vWIMpEiPCWwF/kj02l2B3HvggkACzN3NYhG4qj4jjfq2rtQlklITX
o59Zji9vIlJ11mPVHdy9N1+0MMNFprADd+QDx+GUNEoXHEZtJOfMsq1poxY6s7S9RGJj1qtNHH00
sUOWzMaWbWQmKRzeaLKK+kkVUMdlk5YMK/vgJPBNdrteVArl6vY/k644b+KY1d+yXlb62TV57emX
O0GaQAYyHdBIByJ+evMlyG2HJrygKfNf+WhtNC4eHfya+B/1CAF4IqJi6IgSMbwZGaQiFjQVWeM/
uCZKnUjIkecEcqJz4iy/B9Nlqlh++GmUrKkwycDXVjI2NF6X8tQwzcKBPAOFFiBvXPC5PGVODM33
mGxVb0+ABQ/DxA/Q8A2lkrrz3RMYn1KiCQeOQ5g0viTIOmsixE4+Dyb040UDBuul/g2KN4xti9R3
HllPT27On71FeraY5kDnTx+usN3dyJByFVg9pW8nIY4qPFgdwoZ0kcX6dHkGjs11kGI2zwpqPfCw
rRAy3ZkfppOMLgjvw97UyFtycqK/rM0sogCwUMQnbR/EjH2P6IYjNM0QWP6bDQ0tmFzu6wegbnx5
rFQe5HRGoF49wOJQIetFRPgy3AhJkFWellsHwi4hayh84+oGsrNl5AB4avHmnQTiPxngoJiPuy7+
D0fMPt0nsvDPyRirfONKooPk6LbErE5uLz2FPqNGpVlcMynpS/yeic9gFD5fMd39SmqR3NU7Q98s
RGb0PCanogVOYWWBUKXxRsZciwz8gAakJTQ/YgaQhvbEoQDiufCGWPCAa7GkR0sBaZXyZ0m5Fjb/
z5iH9joCyOMjOxssm77iIf42xIqEh9n9TEk602HTb+hF3sNKdPU8eLYZCoNns/rW/38Gp4Uatjxj
96qdfBUDzltTKFeyHuPwyBTxxob7n6Zl42QC+dUV6PCptFkgH4BwH14GbeNu2U9dNDhpFvrhFTUg
oseZeh3V/X21Xt5hlJl7dDY2GpfO5nCDwI9xBEBPmZydo4RhJf/2tsI253CepjIlmzdXJQy79mBp
qHaly6WyUY/YgkJ20XXerJ6tyuUwEqc5F9J7SvU4qlj5bAlqjF+iSIKyfPW0nEF0JrtJxcPeZ5qL
LmmlGsscC8tQy62Nzl4dw3DuLVwxcUAvUFCxsjhDuAFTClawnKrmS4ouw/u/cD1Krg6CeYOh60DW
mWWaDH/yRPma4UNIbXOB31Nj/1HNSO+77Ixq5zdLuXna8UVbcfE8UFtDgxzuS4tntZEAGR6kcCZ7
Xr+2WxWALgOaNW78Vm0EiBcv4NlQRr2g87fhutVH+mQ/sE4I6kwW8RsUGflFQka413xzOAnn9c8m
Uz7M55BbsZUzGpf6RScIDsyXxxhyGmDCYjjom6JwcIXQ+1sapJijzbz4NLbySLVk7o2We1RevYVR
all7r1l1Tn0WtRgZRcIOFr+KqoVlwEJRyRBrOVObPJb2EObvwSAzBjiWvLaIK3NiQ8jD3nHSztK6
1USxZbjF4Pg6GVguYKs+2fhL0aH9jMUb3HOvSUKhE686TqGZF/SK3jhBQsck/MEpr1BOFE3DM+P4
qkvSSZFPS4LavD9D6SWZyPX2Mm/dbBXMhdiTp/zRal9/1Due3G0WNEDZs/UwNoXi0Q4Pp67+91s7
rEri7viXvLFsJe3iX15HntjGW3UfcqmBLFBh2xo8AXq2iuTF0EBBW/1n9Kh8e7kerHfLWMLBLnO0
LnSuxhozA8V7Q/+H7clPAf7DY9zXDp/KVIc/ZWJ08g6bHNhp86sFkOLwVOSgyjKuYfMQ1nfJfHY4
Xr+lErvQciI5mAVEJyNXjxCOMVQk8wRUGUFlftBOF3DCfOHlYd0dYSq3rEEVCP1nHXuhryDDgaC7
xR5o29pzvpxdj73Kxpd05ZiKmM+mq41eIkikaaGndlgP3ggR4KcuM+eJB9EPJLeth9UftrIwfde+
GbPizlSAbUkAGJzq1FJZ3RFrXKl8RqJDy6X2KuHdwxJVoY6Z6S7sS8i1ij4BzOdHOYj/tulCj8qV
XOOlz9hcGgZAR9hYOnnmWi2c8NE6uWIW8X3HpH7No18VLJblKUJ42IB1U9bcUr6i5XsWRGIKaHMS
pqZptxKUrh2jbX8XU2nvAhBDR2Gzh5LZ5qNNlaNFoU0AAEykoVs//gMmNtCu9/RJvKjy+yeoum9z
DylptdnrumGkYmZP7bk3t9gtDq29eGhD6AsU1lyEW8ujIie7T76NwOSveeJVumyVnEQvPHhHeDtA
D+uz5yKMl/q9nWxLmYGFw/Z49MFZs2UPCA2iqqpaR2U47f1R20HKVhAVQKg2Kyy8r0WMx0eh2M0V
LDihl2wYQ90eA+j1Rx+GLURDsQyEHuYJ3Ncv8ae7zDSdLejbSLGllHykOYT8NbjZGIOBrsgh0pqL
w3hiMQJxn0oxAEUhCfcdakpIplk+6ir74HHZcdBcNQv/Wta58YMu64JjVkEMhuuf0gSV8VqaDwRr
62JtwrijvOBObFBwmzDQWq+9gD7Sigw1/eKJEkhZgbDFh4HpD5HoW66D4v11T7z7Vf1YWMPHgi4Q
8zPsL29fHR10cOekY8sAsrSdBqE85NGK2QD4lH0jhj+2+h9WTZzo3yx9Blfl/YVWc1qYuAjcwXIy
HnRRfUuxn28qJOB+Jtx/qWp0hiE4TxYf60BX9kdI54DpP1Pt+96B14e+p2Q7LQjpzU2DEh4wZkwR
kUtVe8VUBVeT1DVJYZfl0UY90IdR5CJtT2mlZfhCHr/HerSETh0d3YYyjjcTroiOWHgJeWL9cjhY
kunpTHEnM4xucseC0QuKQwb/Qv9O2goQ95Ij7vBRVhG71HIu3h3gVeM6XF3KthoWMMMoKkhqTeSU
/KMH6/8nnDvTSrQQhwemsYEbiGQ6SVfk3bOTVkUKzgcQyp5WcR0L5S1F+jgrzyFtTlVDvHjL1PLn
tAd45X4QsEoB+GyvVK+dHn8I6NHjEG/K3qxkrOYFGCeK+toxFol/F3kX5jS2BiRayTc6sgLyG6cQ
dYo40s/oyNHjeuolQIDP+VQosnOiyU0KQPBBjjQ9kHgzp9S6V8fyWLv5VNbgRS0Zb6dau6x1uavc
sZzltcP8RCqwUlIBCKVdhd2Gd64g5kwwvsrgdpcIob4MIDYlh00CBaU+Ma461uzPZ3+RIPXeOQPm
tao0mbGl9lqNtxBK9nDrhyB3/VNLaZn60mwlyzU3RZM96MPfIrtluSyca3nc6f58TIDXjGks2Lxs
vIdARMBWBEY/DxfzlTZWcDFQIKsRj5r07QGeoM2X23ySnq8N4orek9kw+kR2Mj0iQhLBK2p28vf5
YRiHTgxixg5ympJVENZQpztr4R9q65rEXXro1d+/NRU22qEmk2KXPKxWivLlG8b4Li7JpCQvjnA8
Mg6Obd3CdDAksdybMCuwI/jJxMAnDNtmQ4Z5JJzoWPIfBkZUF3y+IqRHptZwzmDwFyfyf8VUVTU7
1mb5k5iUNHhMvYOU2YAgfwlek6VXrNL0PkL5hEMas0H0e03HoEgUwSDBJCs15Udtao0a+R4hbxhx
b9ojpwSb4fw7mPq5/9xc2uaAkQURk3CQ0GyNVguIOZSItsH6bWjSSqdiCdgdMB+U4suUoHae3evT
IteQ0PvknI62lJfBXolXB0QXQmq0UtnQaJh5hlXhhkqB80iKQCz/Kf8ZWZjERIFN+f1jO7cQzDdv
a1e4i0m9cnj0AtBR+buMmQ52iRCcAF5eKc+hHw8jdJvR7Erw2UsWdRnP4JtH5huscQOQLmpmND7T
MP74/Ib7UZ7fO6S7boNwvCE7w6jDpOODUlDZ1v/uXyyTOMLelCvCRFVDNE1i0M+TMxEvHsQRfXhb
oKCHDGfAzt90yA/W/wbJjo5wdi8jD9kD2SABPVPExU4wSrk9juLEURHzHQre4HM9HrkZeE+JCbtC
tSb95E7wTssjP6zY6W1pxFMDB3ec+IaWyCYD11y6CDAn46Cqx+Evcnxnt/d/xe7SoWqnxAASb5ym
lUbO2Hy0SfM1ghSigAKn797vQAJLeI3+qrPYiofsOHwoaXChtwPTDi1Ipjq/Wz/8/QjwzQj/JIVk
9/MUiYsYByWwrKY3nRufQ7jOSdCVC8O4+3Mrh4A58z1EGkdg+i5VfLaUTw9XymiLE3DKdtMnXVLk
xIbYIDMJJtZkpxvhjH25h+V3NCTnD3GkUDqL8drBya4cGkYTUUZURjlUDRG4NkB6hYakZZXd4hig
as6ib5b3eSW3Im1wHy0PEsG7yW2lXGk/yQ63s5JepBhjqadKMZPc5MqhMmSpPGvnGs57/935zYcU
bNiFKlgltqh3EtI1zPFLjPReU0p+3owaQwUgA03Wrq4L3588ocBwBn71lsjJJH4FuC/T0CRhcQTF
CwvTbUaMG2P2wci2+6QjckcokEuZt8MSa5K4lLeMyJW7wEfw4MZct+ToHAbCYRgF79N3+iVqmIfW
MjZWSfzVI58WutSLBtq2x4L/4C+JQoouW+4usvpn5sPUIisqte5zDkrvI2hf8IUcryYnJbeV2sb3
azfSC0n9PCGVG5aPDev2Q/fjs2VTQ7z9r9ABoa4SMviRHlC3gYjgGpixGer8YGCpYxaZTEU+mB5K
l846NDbJphWT80J9rtDrMtwp9yefQZ6P59OfwM8NIlfhSKjxQt6bTfxIns7DA8tWeGa+bIsMdogA
2Nerb2/IGbvaIG8lfCRBLxcDQKgLhCm0WpEBhAgOfopvrczmRl9Jdz7bHDAmxPOPSytFVFQ3byGP
aD6me25lVCbJF7J9jXmgY53HDDtv4pIUppsoPr/xG/bQe0ePve3Z1s5UAAFaKYJQaYXof+snuvjt
o3VI4wVNR+DURB2TlGN00JtRwKivWsDmQ0jLLNKTWf3q0hbChIkNXW+bPS6/l46K8rkiiYiZTlOf
bY5btYCDpk6hCIlLQRrotLNtIUYtaoHHT2HbvjuR5Nmia1tJjNU0RINwbnt/CA0jGbnvtrqFj/Dk
wpeNbpKL1PdqSWaycthFQwiw3cxAiYN0nm9F71xZTH06CDhkaJ94UOMbfCRE4oveSueFU5mhkfYH
sNwBjSQoK/I4QZHANbu6o9+hDKSHg5w4YvN4n50/SQ3vea8pkB1fpMmrMDSPrLCdxWoOmyK6T4/7
CXrKJ5rp/gzylymfgpvMmTfZtXYvcjN6M85FEtO1wbtxpIVfM5yml3sfEWjCWHdTGqt3kyjk6z3Y
LyGIGLt6LNLa5PHBSSvKlvDTUfQuO+vCafhr8m3txKJecXOE1fP9EcAg5uwG20F2v0xrrKYHr5FR
TDbhWuaMGpvql7gAMMnpqJ0bwIVP79LzpveymXIndATvDll/rNpu5Q27OZsD2jClKVmEKtmTqlH7
kHp6pUcHkEPbvg7zmoXvqS80Uuc3kCdaIWjoqK25wtzc8r0Dbx+E7GcTgfi8qKWfSG3q33Yk+3kD
O38Xc7SVGTL3KuL+Tx/bISYWfhGfXFSr0lkmuZj/rtXVDL6zKpV/3ApOHK7SdWi0BwyBzAfxSWVr
zY3R5fdNFsAPH9gXINFQd56KA2c9IZq30A7xmUyHYol/hErg6mN5ghm0dXky1jBNRqYAVCQ8DpJB
pYE/xHpYmGuKJLHGKvQux9VsiBPRtlvUZVDwGfWV0gJyzm2Dt9lRPvadaoRXHq91HDh9swAgR/fE
8u7Ax7pOF1feSpk993r2+s9DivXnMGdOoxxJhbQ6AL9ASCDes3bUeDWnr/uungFxi9JghGYanjZZ
zy8t1fsG0+E28lJIYroK0MQMfSEKNvMi4HI9O8lGd3n9G7gOn/FQZ8TSOJnEpRJzUOQU8JgQxuwE
mjyHhXolR5hhwF8KgDTMVREZBWH56Af/JHRJR9kP3AS5qHIM1H1Mn0Kte0/F6xTT5vHllsGW9FiV
FWlHYRf64QRW9yIdldrMfy8YBqc9lsuWQxcUiTEC3yXeF9BqMlkfJOU/phATv6MOB3z0Ok0q6PMr
HWd37QQlVnmcY4Kpb77RDK8dGAsXWhDnPw61HGCqIn/687FAt6xL+NfcHMFdQfIlZTktZ0POblBw
tGRXDYXqhqZEd9J3nwBoglWvDZZWtaPRvJWcmYbUADx/0YaQ9xP6z9A8eNSxUElesfjSExTDll0B
uC7Jrab/mSOJ5CGTTq4YM66X8s0JhMM8pxG3112QrFWbtFWD+BrvYurahqcpJ7WRJuvwb6LkNo7h
3LzSSK92lZcWnULX/VEPW+JFcjsmZL5QIlK+5M+ig9AkP7dwhBISLjAzX1sINxPY/oLXEkIWihli
Puk29c/XQCKxFM7BevhhUaq0t62AQaCsYe7EBQGuo6UFFxbdFHKK0z0dOq5sJNcz9c/H/E+zSzbq
4grcgbIdtqTiZtUCY4wpdIndLPJwwdoAr6W41zbQvOQ+1wDOAHeyi4DupOfHTYTDrNBr9SfznncN
J9PIZvqxCwgS1DMAgqiP2U1gVbFsuKEEIudvIi9vCnxwkhdCTgjbQ3OXfUFDaOSixdTShD+E2GTC
nIcFhAYONBWhN/PhHTJFfceL+caTU/mkls8dmBZM7dmzxbh/ee8uj/KMixTLLOWZAiQUMx10ixe1
lL6B/O+b8Es12gnOwwP6uCfOr9Q5/k9CbsHHLqmUrzespn4yCG5Yl5w0YDgtT8q8rZagHJlW9ZVL
mzef4CsKx12sUcwZKqCFB6Nc7pXDJKfYbxnJONshKY4dB9gN2cqKvLYe4jXJ1owIV6cwm6HS8apV
FTyiEOxhVIeuIr0FS8QH42mgrsNsU2514vQ8f6xJrlHxtoRQyDJdrWfuPt045xHWIjQ0Ba+mx5sF
S6JMjEkwEYHrxq9dwtb1kuO9VtlnvAm+uQeLIgA8tY1cOTubZEdwVilez6x6MDdUquRAHpWRbU0V
QKXXuwuAAVa8hcGaCFKQYpFkG1D4JfkzMfZjKOr8Of63bjzxR3exVcO7Avw0hJ7IvO3Nv4yr/5Ha
JxeNNhZIUCdE1w7L770WU8Pty1vdSVLF/hKYyfEuJlhR45VCLTIYjIl3DiXTrUKP4O2Fb8MlpB+t
T5hgi3zmQG0GPU2qPIKNdOk37TvGLMSpHsZSaQD7INFWvlYfxddaMZI2/bnYVrKpxOctllyRzaFg
e1bDdtKMEB7iAcb74mwSnHoK3TPryUGFNDmK8O9QlLCfUY4b6qmJ/z3IBLbiSt8ZsYKDKUnQHCfk
bS+kwjbQ9oXbZAdKTCrfD7ug0Xwf2YUuyCfikjFN63acCsqx9gseGhKr6prkXUox/EpieTuMGwrV
GE7BAG4Zw7GD2tadHotmbC8P3VoW8lD+T/yR2QjsRBnZLzUMQYxBshh/LvwzsvBH2HzErve+bB4T
byPzq0HMEknIx9Jm6FPX/griQ8J4nD9uAISZiP+03ka/Bac1famImZSAYHWfsrh9ivysPbF2/Pe3
n9wCr4nRXwTHVFgu2jwb6FvUAaZsOpkdki3yoAOx8pOZ+8x9itNeHV5Z3IaN9O6Af79a/YqdZ2cd
0PaS9CjuCefKV98EUSTriEyp5kdzFjK9H7LDt9qj8V63CoDRpJIc4BBTLTC3pJDxxGjTHrLAJoNc
L0EozanPB+DKV+in2GonXOA5lKL9esNVhLlBPgy+1iVW+NloDVgslV7EBWpF2TNDNN95TFj0IOlw
4fJnA5d0mdqDGVZQce10rN7Gy7UKF5tQgG3WIHuTfTEKEnEpNlAkrYt5Z1LN4VYQi3GkBVhr5wEY
ex6QIhV3CMy547C6LvbIxL+UzJTTHVdggaiXcuC0otuXcLByP6X4pa/xacClXDFhNVgaDaZpDIHO
vvU4m+h0s2PWFRPqJOX/45PZmnuV2jMjHiTlTNOVBPjksUINYbh4XZiqjRxl84faZCwlj2Lh/l8/
P5arSDK7mD+AycXpWj5Y2y8uXrfaqSTN/hOFrrf7EmnOqV1Aa8NMf5OAEldZqjAE9T8ufc9SM/lL
KNMJdsoDfe1pxMxBI26RPXsXEi9hxdrndsY4EExisbuBVVUrdNmegJEFbFcrIPrUnV5TCew098Sj
HcATmI9hVYBL6wIV0TSqHHFYW1pQfWtnfL833LDR1BjOiIof3fVfGVroafpLH9Qpieh3oEckZuFm
hrL5O9+oQzwgEVtx3UcUhBxTfHAxdc+D87iXROuPBrkCASF8Cc+2jy51HzOvSKG8K7WHQ+s2T343
iPiLqZZhnOcE2yPw+isNr/ZTrzMzUz2WbqZhaXgEcNkA/IHRhHynCJtfv9cKDfFgxeJoozw7Wpfu
CcIM5/YZUk615hIP+AS+jcCdZhLTrH8Qdfr5v4gvxpA0WI9liSg6xqYfIet2hboMfE093oMQ4BMd
5h/uaVNTKQIHQx9bgfWbDAzbWjbh3WE5qh63m2KFslfQ2wrc8gc3/YzaPLCXmQVyS5N7kpttTkAs
Q2/fSAE67xVtJi9PSWNhBu1JCZGB/eEsv0QBYd/zzctrJix564kVvCPJ1xoe8Wk9WhEXGP3X6Fpl
76nrXkfyW2Pv0EHU2Imrd55AIB6NPYMExA11cf8AgDh+rO4MIChrCGSdD8FRsC3RFTrzBsjy6J/w
ovxnrOGHFU8JUSUqP70kIZNb141N7CrpT1hgRSqwxVbJ5u5yB0u+mZ6qCZXVfufAzmtznCqmzhMx
zK7nootVHunNH7ZPTBylzoEqtV69YZfU/tEwaHZbJgaHOgSjRFyv3LABVOiKLv1ygMgZZ/V1oGNV
6LCWqq840MR+Ldsx4Hb950hSSgZj41ntGxKTusr/onRy6pQyEH97YefL+hpYczUCwBX5G8RBTMZE
lkmCHRUCIITFmIB5BMruwz7SoETJ5OJQyjoQLWDXRYS7OEmCfrgS6jb8ToRVmqtz1QRvX1csMXso
GfkqBg7R8Ou1tZxlO15lSgmapc1Fq1cM6FibHTl+1y5rfyO6N9NlwxtznpryTKtYSiWyAgACYN2+
JSChpfIIxG/cP6tBEDlFDesE+MlzbVBIs/hEI9kILMVE6v33Z/R6IKQIlw0kEGpmfUmIiwftKF+8
u7fxTxapDkFhddtnTNeXSgf9vgBn5XSyuNPmra9PAAxHljeiHjhXqmzrBwBSoO8Psn2D3b3L1+3e
E55dVD9iIuKVYROP/ydb9OHrfu1NZ3m0+ltD9wBbCYwSlTc0OgWzBZKbYss7UXBLpgv1pXrsx9fq
0jQAH6j6WsCJMPClLwh773KV13VrQIvHPSXJ8FLWbXOGYVQ1km0CLJXgQC6VZlGbNrv++mHEpH+h
o3TvFpomkdFVmGEi71cWxP3kJaCpwNcDBQ4pgpUuZzPMLn+W1kPhZXHzrrzCzce7hgq3CAg54O/n
zmmguKjsC7lOdaKKaqojGEPpC2wtKnBNeGsIRJwz91RkID1qRGtB5BQ9UdwquMfH32j2dQtCuGVi
dfMlI5lYNYwhDwoGDgRXxq67B6+2Lc8w8MimeXkxPS4ohRW4HW3lJgwvw32CxjDe4q9EpIyVCF4T
VEhPYOzvu7R+bz28tTbvw5hmn+lMAQS5N/Ij20D4krZsnv+e7MJGjlrZ9T02GeucUqJa40D59NUF
TG7rt6nYsbbM46ffvWRXbBh5oHfG5/06rfIx7GibIVHSY1BD0/NfItAb1+euvrhFIQqiU1gJ+hPb
Hzk9Y7aN/7RAyaw1ARrbXwB4yB/5XxKC1w/r1REXJY4RMnxyP+Za3YNQdsBEVbDI8ub6PbCQtYJW
FPfM5TpUCGedWmhWVk6v8RlB7fGWvUkBibEJI6B+VMvP2Tv1LvOaM3glBOpynBADwpfWPLsgIwTQ
oyEBqzouYE6KDOWRl0uowv5i/QCqw6QUJ18cyb/XwhFub/pxpZUQ0AZysoDFtE50cIZKjSjQeTmn
T5uHcsMBRUs1oUON3Jrop/+PIgWXy30COAc0KZThCTwSgnvLVtlTF/gxij8yAOBnmE2vcS0Z43fG
apQ2F8zkGwn3NNOPSeRMafH9xQ5WEqUcKrdwgNGeA5zEhsAdMmQkm25CAV7aSIq7/vIa1v0T5vUp
zVsIFPCMe8CuvshVc3xbNXmwNoFjBS+8eecj/6tZ/Z0QeaLUeDWxX3fPm1S5TaStz87ff5O8W6g9
I5OedO3rioBzvbNiX2zFDQ5aOq7hp22ibQXDLwinz6g13jMv6UCLT/B7B9MS8AX5BvYtghol4YfR
KLrDJDi2WMpyDswSWopAKGKGJhNfvBNuTVh7eA97rj/0tEOuoas61IHdv470Rykl8F+fLbL21ZXQ
fch1Zzz6v9+FHFsqHx0Ki7oK+3YoylCUlR7ZY4L6irqKWmyW1iqa+DlWzaRGBBviPHkUNDUptx14
UpwP4/HSNR4qFU/2qPT/I0ADidb/Sq0Jf3J0FsQtF0iaps66OUEHWEaxCcCHZwFCpktMB+mw2eV6
1Yu0KyJE9oynROJVHXA0l9HxmS+Mm0cG4tN7QUSw9n9d6UHzdTY6JQwtS6Atv8jLRrVW5j9Lxrro
LTazBrOgg9FJg0E9te58GoSMbcbJ6Dvr5Rg6H3F6JbQiML6QCYErV3FLgtt0Q7QS5J2gkOAa+/qe
RphYhC/6QRqKq7RCu8B8BrqDCqgWxIdKHlYiZQwERKR5NJgWLS1GUaUQnhzVY123igEPMyNGfYpD
TW67ha0cqQ02NOEQZwouc/CS+S1jCLM19K/jQr4jB0OTNsVFutp+qz/GzCu4QqbzEDoK96nkir+W
NZXhNIhj3i3b2rDbrVANmtCedWLcHAkOhfRazDyLU3uNWAf2UN+jsCRAoo21Bza/htdpf1qB1CgF
K9bqBAVD2QgP3f2TL8Bqm12VtSVqtviEcXOXRx4CC4CNdG6ANztlddi1aGjGit5wDXj8A/a+YV5u
kMlupQIrJ4DLld8ZoB0z318bMk36siC79F9il/MRob7hf67jzP0x3zdxyUw3lgCO0be2SvwoeYiV
Cm10zV8pwdCH7dm/6PRqSgcRJtfz/vnw/oQDdYzBVLcnE4ltnaGIJY4pfA/wKy1T2eZsHgwZY9gF
pMCTNVw8HkyXcWc6nvEHWiRYcrR9YRkiHCF85P6T++8ERerPWlQ1r5D69o7c1/K0myc09uG3Bm8Z
QVgWmefbjLrs3mYmr0HZv2vP3S0KtlXf2dv1ZLAv+qmZThtX78B5UwRgOklLwkqxq0WLyq0heOxO
50yVCsCztGDfvf788AiUhCm/yQzUIwOmLl7uy+XekD5T042ZEXqTjBiy06YmbZKF0+1chH3ewL7+
MS9m0a/FDyG+n49a4MbOdnLWu9H/sChzupDIqHQ7Hl1n9yM+9CNzSDpBM74V/EOOuR3hOwoPE4Je
buvheqzceghVLbF0Ml+B8F0xez+/RgvGEvjV6BV1HNPAVZAnKccwToJfHa7iA5uaCnqsl4ZGVmqR
UQLpMVz3jScsH5Uvjp1okdDQGOv16ks2FoTXojHoghZsv1gNPnFEOJGycxe4mgWAuu5En98kekoP
744WlwPQ/gttfK8sMenbBDvEYuQprg2oIzfST2b+uOdXKOTkJK24xLrfHFzQAWj0F4/vfLLca4E3
vVIec6uk/d8oyIYs0QltC7Ea3BibWADX9Wa6SMAKOj3PUnG5Zag0Zdt84nQHkQmJIfl6Q3jb31/8
xqWrAbApjKSvPxnaAequww2OWggOU4JllWA6ywKmp/q080pNj0Z29KCR8Eh4e0N2Eu87ycLQW95o
1ooGzpWm8MiYVirF3SA0RF8y1y2MY4NNf7gT/wttKW0NPPCWC/H2KtYC+yYMDvFA3wrO3wqy4t9v
pKwY36c1lBrU5NsQSvbfC2jVRACRry56tw3aJNwFYJjRYnJ5L6Xo8V+NIbv0U1HtEUEg18Lg4Ox1
r1w95uQn303o41aN31VRKgu2lJLQ4rCHRV7mknhphe7QLUg/Bigeuwb42jp7UCFWdQynIkTQz1cu
RAbnvC7HzC//fmSF34pdtODl+sat+c4iLNNH34htfuL4FDie4xNbHiRbg0pTZSMGRd0H/o0nvTBM
j29TqWKb8GOgA89LMroU4Qp59XQOPR9jR6BPNMmqun3ksuMh7AWfT4DrsT1WZIL0cRxpYL1fiW89
icXcjbHzV1ecm3Sf+GW5Z3OlJaBEuMBB3iR8rrGpjjdF8kdAc3arVzEECO+KysJaLzIay8E27FUD
IVD00CUTxOhoCkSGq1hm/oMvtLJUVgDFq8JXlQgzEeK/eQScq6ad6sPpKXj7BjMVdCCo/X5JZ9Kh
EO94aZbRnpCUUOthkI+YIjzOnJ20+bi6Ast/alyjytEbN0sX+aBMUV9pa/W43+mvY2xfiaHL70ej
aHfQu9j0Yt8iV9M35J2C1r+r0KEefOWiEJBECYXYVbW2KMMZrUCpEDcz/sMsla79YtXwD6w5on4p
PH+IunsJ9U80cata1Mlgfkv/Zx7kA6lMVOB0+Wb2eMJNYPRhIPBwgZTqlxxhzssXh/BfSd0hoU9B
Y2yND2r0F6ijwyzTsrK5zuNSJ5jDHMxT4gMpmnn87bHM7giU+ZTPp0xhQAKYZkrZ5okTxwlqArK5
GX0hugdaVYdBT/gH14WY6OV/9/Oeip5WvReJDgmiNzSBgm53Q3I7io5m37ZxJ6AdEHuyGJtXcpat
q5gH+BroYX0He8sc9pnWkenscHr9M2b5sn1Vo/5/nqh5qUsb1zOw0COtv85ssCeMcSmG1VtYie+3
Tlf9SnDrd0vt1fibX2tN9bRwzoTJQHS31TZAWmAScMEFXiXUNpoMDaLnO7NjiRGUSGk7ANsrSkCh
3EsgIL478TYwVqHNCERT1qkB9t//UWrOdhxykyP4AEVw2OKgLw0GQHQ6nWclzKSXSKrf2GeetjNj
Z5le7UddwhgRwpnxMEhpsaC7zhPRbP2PWTJY0r5AlxoBFqSuaNkEHKh7E+woq4gLAjKa0FJKP4C6
nfHCzwjn5QoQBwnV4Mc9G351dovBE0dFf7DEe0L8pEKVaKj0XttrLUK1EEMyoaueJoFVtSETwO2I
iCtk3R9ki4tQQxQn5uQSzujJ4tVDgP5JnYGpIPYIcNdgLEQ8wG6lmrovmHUIvDP37mhZxcmbbVyi
1z6ZgEnADlpyiLUrrxJ2MrmbYk3lE8k3v8r4gLPv5Hu9zUMp4zSVCEQqwjZVPVN0TybJ+asqZHlx
mUKF+/cKVx/gYsOZ+GXt9Ax65dCiwSVzC5q8dn/TIVFxE5yweuIZNSZ79s46nhoQszoSNnERSULa
PpZu4J8E4BJEjSa20Ez07VSx0i0dSzbazAeeXx+vyXf2TXiavihb4CE1RSaHfihnHnuT5ZrBNIku
0i9k0oH7kl+3yPCE9Llx7/9n4gKb7gGhb1f05PpdtBmUvQGRbTGQr/wVOLyWJE9LWxJ3gussZDNC
20oEefxrWC4kw0xHIRD8RM+LalgpQqOt/loDRl6OYyAnEeS8GKeWJZu2i8wPHujO7CvxR0SriUkf
myS8q9WmPktXo2JZMjFt/uTXjIDKc4l1a3SfQW8gx+069I4ZfT3VsHZANyK1dNqayKaDB9qReyOB
Amdo37GyMk656BUep4TbAXw+tE9cfDkcyMrqRpMlOSBPp3iYri6BSSKrq3P1xfzaxpQiswIEEjK3
Bf6fd9NI/DggnPLHU1fqrv/orNXEeZVkzdoDlEZkiqwieCNnggykDeAr1AYlCwmu9RDKzUhx8g3r
gnShCRhARFDwzBfC1WpTvASudT3DeNsf5yZQwv7wZYTwCpJWuoXJrlMAqdP7zVM9/EhiWBFymCj3
n042ZKB9b7gm9AG8CS4waYbJj+ejKPkvXMG8pG63buJN1OBwgkwqTwkMd85n4jMSyG1Lvqnp/y+k
uRvGkM3iHDLiU8MzYWChlm/LyymJLQ2SbMbNbyuU13V3nwyIsM+YZwu4QzvKHPoPEBZxd2KwrUb3
DjwZxp3+1JGJr5VaoyQWZxiU4a+72A6obcBFNeUp2ZUObTuZXRRS5f4vilHMMh7M4GmEXixqT3p6
cz4EkVwWavEdPfW6GBDzj+TBzd4LN0vrdqhjeCvECdGckvU8UnZd7HCBno1poCxvXNvZoQ1r5O1M
xBpGTrTAHqTLxB3c0QrpJ4RpONqox5lKFJgoAxNi6fciFCcM0s+dYoG4B2MYu18ytSnh7U0lW1r8
49WPy8DlLBnG1O3Mwh0XFZHAuqqYSV99f2NQhsKqmytRuTg0QeNgfb16E62h1H/1+r4XPUpyogtz
P6RMt9EmeFSRhhIdBRUmEIJc8gCc8ekEOd61VPi5a/9g5TvPiRpuI+6flHN8fZ8ghFKIDnmKRYLD
omJ1g7i0Sej13cTWD6qzkUc3DyEFSkGv1w6Kk8LvHd3ZuOTzagir8QMpzLVkQJTmAbew8oYA7UWC
8tRFbaZXwFs1fYpArTjmAqOL4i4vZ5fHsTCwZtrEIfiwbMhxHEtZK7wDjhQxenwXOrMlq88zkTRg
ztgRpa/mcszRy9s5rui77lF97BhOYSPIZ7x2fQUc67N31b7lc2iczvSxn2zO+G7WkUvr8Hm3CQeJ
ibP8U6peFTWVc3sI8ATsMg07aFwUPN72pEC49GeqlO8kJt1oDHF2LIdW/olaGPu9T7xaFzeDMzNP
jpyCj1uFhQVt2WysOl5ovN1tRiXUzQq4R6IkdDbygNAbQsDJIqMcGcfoT9r9sbXm3sbRjo+yYSKW
pGyJMxRJux7ItJpQVdr+7hrjfdrzrFPBbmrH7KnFqmz1SMxku56fe9VKJpKujyFz1npPDUkIFApK
ZB7NiwWvaGU3aTLXQs463l1e2YRuZc/fFBmsa8cDEzR1DXdvfMRRM25SxjwyZlQqtXqppOVO9Bpf
t5Yx2pcs0O8hkH0ed5NF+NrbI9VB0vTO2QI/JF3vo3oF6kucs8JAK+V1n1P1ywPt3Q1DnKyLw+WG
XUWzQ6rga594+I3NgJddqThQSK+TMWOqlqjyqFJRr+IGuUV009b1poF1/Skmh9BRm+opQFwIs8Qv
NZjscVcASgAyk22ExTs9GoEMPZafGcg2KXRfIFSWeggYUM9sQqS9PLHeKGsAgqXG0wIjadzwJOWM
aaBmBAxMTX2xcaKPldvx4WfScrXUJoG4old6WmagxsFZa7eBd1YGvvCGs5YY8dn1Ex9kG/M7HVTy
vUfkWznFGRFAO98xHyN9rzB2Vu3mlzN6EYlUO7KgMh41O0tn8wn/WzEw+6/YZQJZXFL1MZPGusAr
bo0smtt5YQhzncOvCy6KzgTbv2D1SkPvHuDQIaK/FjsyAc35bx6M3CNEQlFiTCXWwneWLBoyX/z/
+DpyYh38zTViM9Bf7VdcbQXzpwpJrIkK1lgksZC3191CGl57OZceTJ7So/aqPXZ5s0qDk0sxYu12
5nlCVz5hgBOcixw9VENHwcz/D49WQqHFx4tI2Q1TGdoryNfVT607Tg/YpldY1bWZcxHKSz9pGwAL
0ZxElRBJq66R5IQhElkN/WYie4vO8vOebtzM5jp2oBgNE1OYl+RUq5GFbVdqRn2anIX/6HN7/d62
aasj4+NeKexyGbL0Qnw/u6d4xILnF+GGNBhShG9EIPoSfj9xN/BhFPdUt+q8k36kDR9oDGGx/Vy7
yPP0yKYlwTHtyZMvb23YefHVMiFOCxZVXPc16FMMpW6+cxbwQEY8wNUY6oczPxgpZT5sdyYLoYa5
pKzeCjLrKNxHY2MAVayxvdPsvyZEmaOIaXQOfIcKWgPbXk8O0TuiWOfwtEMwGjvKCtobY1lNHXdD
+Ki1MkWo5VRXVYt0heiz36b2xJitO6s2xKC0lDnkMC4KoyO1SDsVT94shdmzMQQ/J7yaWuccKao7
E0CRUqlmQpCalsHeYabWEdqSQ0Z+85WVB/9CaDQbOall6/CsDNwtUh9dWlqMBX30zAJDvtdcZE/K
/KA8sDTfwlL4pbmMUHu7EV7Kye5vt1B+D1CUcUJQ/e4/HR+e1sx4d7SXTLkVZcNsfM62OSgkb9Ly
CGG6pTiMrx3EfvddVop27HJZ+CO8sSEwOocGsXxbSxb/3GTLt96wI4VYVSuTUFKoCgjlrNAwK5sa
CLxTs00sdwZzFO0bueJ8oGlJ4AhhJSxy4n0kRZWnCB3gHzlpkr63CiqaYjIGqYYxvZhme51kADsj
MRmJ7IVuqeMk3KioQzxeZi6LJvVzSZnQI5awj1+PgosAPhdbBWz29fXaGcAnsXEMWQc82TCnkDoj
MH8YGAJaXVdWqsISvJj9FH+C+ozJWpHdutGdG3hPx9awa5Cs2naVZQNZ5bH+ySU1K4yGNPyGCW0P
sCVEDnKF2u8lPtMDa/XfzjaGjfLcRlq7H7rWppZZK8GA9lllsjQhpuorwAf7ejv+Mo3yj+hc+3TX
j5sedRnNNqGNQfH1bp3WBe44fd86nuGyHZ3DoqOmy/OJu1bDpQBsD3mbQ1NNqSdXe29m4FqPctef
eyiF0LPhRYjhHCDto0+wDzTeSxdpMJlgq27UE4JXKWcwrMzg3EOw9dBf/jxcVLGqTxlH8Q9HOmT5
+emQ74XI+g3/SSG4AJwBCA9dwxgV/V3O+OVaAEBeK1HgpKw4550K6vV8Y6Jnm42p9d0Q2Tr5rKu7
TbwubBescMKQlRAelWbVvF3mpDN2TsLQfor3y93NNQuVn70n2Quf7WBFc/Gt/K6Id8KjAQQLfBQ4
keH3/A/Av5KbRgik4zCFcho9IsAIfiMJVzGsUX/2ZtyQ6GkEF8Dh8nTKWbnny7MA/DrHtStgAVTX
JyMpBeMyoV0siYAKj+1fQUREkV3SEm/tuO/GglhLP2/EVFxdHD7B8VK6+HgE0q96884aZAsaZUNp
CxN8zn9Z/C7OINfW/639FwKdZjFY2fPMyXe00Y5k5ni+WZOu9kvfs5T8g8D4pKgtujtLAfUoymSa
D0iKVaWSMuvsybBAkFnWJCeyeWTc68WnB4QM2KTesmbMsDMvbUiG6nvl+lkdctCDTQ1T/SDKrR7S
wYCYBaYgN+WTjm+xEu0OiVYsKbAIskdOoD7/EigKeD/dq4mDw3Scg98mewlOcpRCpMBMNzpzdhV5
Y0p5Vmsi3zdSdCbCEXIrGucO3+BUFkG6dkqWbWzRHZGZdYlnx4gOKPtCaPLevfwKjqcgU8UBWCQa
M2t+1JXvYUUpR6Nn3Qfkwsbt5rgV0TxwwBgbq5zhv/LUKvttAis3elVyRnp60nM4grTYnZEIOS2h
4cZbgb6jhwhEhXesc0/Q1bZ/d4qy+VzX8S9Hc/1ytOraV/ClvmIrrph0TXaLgdVkwjSZ6Qfq3NsB
Z7hSFKjrlmEj5x8Ai+r6Ji7osUwtPgtj7akT61ojPQUW3STqqERBG67r7C5XB3GAdE9K++kaRkOS
/dD6dEcY3FFRlQjRJ8LC0bv4nRb3M0Yim5x5jJdrAS0ReQDyh8qdt7/Q5dhvheEKaJn8DC9PkKj3
txNB9/4CgDWIhmgI/QTvHyXzFyOIXrauqoKu2sEky/HmJ+ptv0miERJI2NitEKyiUgRSBstrgQzn
Zaaj76+BRVkzRaxyfX/xqe2SknAGjQA/VOiCv5Zvthe3XGJzGw6NamzfQOxNrZdtDAeNXaIElBKu
cezuB8UjQMwv3fF1Fz6pResr+K8fIX2v5LBPyV6TknyaTcVE2RopaiA5zEmt8g72CcA4lJVfIbK6
uq623ujOMyXUXpyFPoiAUL32QtKt7Pbad1t37GhwSCcdP4x6FB+cGUW8qCT/KeMtHg6BVobzh/Ne
8oX+OM1Jh2UHnd3EVU79pdHH/IO4kpWFWAbkrui1ABYi7dcI/GvWeaZ07+BfyV/cGQa8v9pZ8Eod
HNhGxU2OrAup8JYYbv8wZCUL81culK5ZKxNF3H7rM4OtoBVXXbBZwfngCn6mp8D37/nOs6PIfl07
uiJbCtWRCCU1EQUm4iiOKJOFgpLDY8s9EQoEMEYvWaL3svhQDUaWdE5bfZwR0GoSj/hrX5EpCT86
uzBMUC8aDMWA0Cq307TT+PXhYamVU+BeqBi5IkdYdsvkS5TTWFxqTKSPLJ5QcyyJUdX4zzSLoIQ9
RGj4XB10gJIi/rH7E8RdTMoHIEGmJagb72CqE6rb859q6M4DxmPjn3BQU4HwEo5FPJkuGJ3C9hHb
WYLp218Krk+q/DPIxj+mfSNHPQFp0rCKa+xlJ28YMlmZznyt0TDMm82mNTUudkFxsoU5ehr4bj5p
beo1A+83TR+lHpPBx8dfDw8obfDcZk4SbjqlP3kLVRDfuhjqHcEVPEWW6IDclvNlahtQ6493opCy
5DjpkafrepjHMCrF8tBVPqFOLG1zA6TUkL/lD0vhqr5h89e2bNAfer50lkCLQTN3l9qlpYbGOIzB
aIyH+yPz5EwJJCJF3L3Zk/m6SCm9g+YPAC9v6CApYaT3/CC9hh4ckf5k1WsKY0wlbZeEleGMRC+j
qKPGfl9tUOwxJ7JtII2hTCUC+Ol2UoyHi++M+L9HZd/jMhsNzN2wtvbvx9klmH4ntveaYU2SbXQt
WO4zXF5/HsLLiisqFLz29uQ5BdP1s3prDNNpSS/+SmcqABS3tDOLgkgf9TnTE5SPCfYqIBlQ6E+4
hERfQJ6Gnch/NPDg2ZO2D4N08nW8Dm4Az1hCmiXZaaDVBgjPAkBudC5U/3G5vPRWYwZj3tT+K/Fc
5sFWtJtlu6sxNVb4Ax6X4BvtG57zBIZSw04Nk1nj3KRajILw8t4hF1sEn8j3/Tv6MQI0MW1mZdKc
mf6MAHra3bJ+nCcgVF47Hn953Eb4JndEvOSPS19D66bsBG4glrnTjZNPhbZC1kJFMu8tgY7MTGIN
0gnuXmheXEunDWgYWWt5BuLGVDLWer8YqahCeFyHVFfvzwcLhHtR6EUUPIuu+t8igIPvPh6/HxOX
Xl/UUr8G54dRSaMY7mIeIapGF/zm5V0bovtfCKSjdvtCWgdYd4RIooeSn5Pol4kdpW9LIdG6+Z3u
Q4otMqR9w5x9/3GymruFsHZ4/iM3jVAunGs72mmrVzLHhqVdl/L41HNQkVbIZIrAqIZ6CkHfnc0e
LqJDp1e1VjjA468W2uqPLOfuDgNkKY4FH0b/d8r3aE+P6WybgTZ4B8SpqbyyGPAmDrFLQ4tPGDxI
93uvCfRz3FjKvooVM3stTMBBnTyOIMcRzUgUcpSUL2tS6z/iZ3u6KktorMChEgJgxYCiwdfIvim8
He978ey+KMSql+Omdj0HQBBdBPZHApfJyCVqdd+TK5LA2PCtytgiVxh+28YsMVOk+qFF/Sc2gNiZ
LBZcRVOq6JSRU/Pd0s6trM4zZxkdabvOpFD3JLDt9fEl3/YxF0bGfBRlgnZC595cfbWirUFQin3l
GzUtR8YFgGu0a5v1wq9L2pJlFMQFqAOFRPiT+pLpC5dd34z7/CpG4pr5u6aXNNo0yt0KpaMqYqY3
vr+CDd09jrC7WwFMb+SP5G+Cp2Tn7Cz4dW1kSCJN+t07A3y+CPsfoKx6BydILUoynfMK9EoapKdT
2HND2zA1Sp5A5lNcHshk3+Th3stwIBxv+UmzkHF/973VCVy7RCJcq4eXVc+9CyHTB//uNg92qFvI
nexA+kqrR0d25uv2xU+ZSV7aIrZlwSGWNK7LBvINhzlEWLje4O1lzYR1SYQoxdNS7ShD7UsV0WSe
aBZs498edMbkfrBTkHmZ/b4NA5hOs9pkzRHRoyCGLEukXZvZHOkbZT2XZRr/YY6Q54mM7stI3g62
7J0XT6gNZa8n9rCQ5VtZ7VUaRfmiF2e74W7WTp4rpQ7zafpzbUplwQ46y3FmZrPpO54HfIQ80fCY
+NH19E0tNivIZ9ui0LEIb3ivsa2gcsbIZmSgiPBHWXV4YNx7q2FGoP+LOBwQatBJz6VUD4LwLvUd
Ic1I/NDd92uCACYvD7zmwXpFAJoFIS7/9jFNWLoxLmlJNk3u2GFNcUG7er2wooRzcX/eGzETgz4l
n503ccg7oCDEvj6/zPTCWsnFWS28c5VjIjjSqQpMPtnW6pUWVtGZn/Cm4U/nLK7lRV6IbMT8mwey
+kFS+unj4UmNtX3HrxJL/Z3Do3Fywpqjihl6h/8YrCHlGPcIEOMbkNk9DGki1E/Kve7dgTopLrAJ
R+wLt+TJXQQ3eEistcBL+fyxu5RrS1unE4NBpka2ZDtbdkE49FYHbvAaiE/sGk+la4/4h8iqmh8y
B4p3F+j0VYmPQ8YBJcOcQqNcqpKoh7JaLzPnhSvFoDvnVw+RykEzIkWRRMC7A+Vs0MQHDwE8W42/
j+QxchQlOY5LPbpVJYUKruFo2O3nstR/XfONNhJ8MZTA6QdncQS8n5uT5OXZDrcla55Tg0SginFT
Y/9W8n8yfwWIRhLSehe+ePslBXcXvr0GvPtHJqJjZXxYFG6AFMxTwL4KBRkCcARZLTAeh/gOQndy
EA8DlU3agHfKnH2/zpuhb0iHwji7IQ/36ZSbsp5piGJxsdqaj0eOyH9iBKCMALFtNuqkYIAFJTrL
67zI/PmPhffH6W9lgbqtUDZ4XeY1DCCYxf1c+4SC69KvdRMvuflRtk7T3ro0vo42W361+UP2mJ/6
BuzL+Ln4b7n+GTQP+luTeRsVUAE4jNuNJH8S+iqjaUeBjYVz2Rs5tUe2TMo7TtX22l+AAZhHjYt2
lxT7LI+okSoSd4/3suDOWl43RmWG1uePWUDkGwlPTA6g6gxRwogsmfuV4jzlGqqRFet5ORuZIzHF
trKvpJhMNwxoqShRWppYJUAysaiT+xVchhnjmp5ie66lHlfazooZtu2PanF2h9C5gPv2ErPPJMFM
4K6EP0dPveCAfNOwLSh46brfCjuT2ts8kC5ejNOPfZAeH/5KnJ1HbpgGzN5agAM7HIyJe1Wzjs0/
joTagrD4JjR2snxxXbLrb0esxekzZmQyVFS8+BmmEAEb+zAnlXJsPkFeKOly6kPQ9vnUpStIhelB
p2fHbJaqtb4+9jsMWe/a0EnoTzG6BLpcsA/aaNUf/cOVdNPUR8DnBo1lJBSTMKe0lFgoqd301ymM
zJQmi5lKDAhOlLlaJZosOUPOJ6HFaozq6ohHFOOVzGr4mTk/H0mh6uD2F1BzJCpAi0Fa3MGooPvb
39CCrMDLGPAG20mbMJEYIDjcmWpAM6sX0BCFyy8F1hXvkRLNHYShHgoQdfIMqh5oyJc2oEIiS3uA
Yn76C9M43eqkYXtZqo12R2aFLrQeYn94ykly+hCnDc8NZAC6McmXDA6YjJR5p0VMGaKTXxQn2bBr
5ARzQwHnYql1K64CkX0gBflgrpWR6CK0j+VgpDd7zFbBmwd9cgBm7OuAyVQ+ohkq4PjmpUaaxpOi
BCZEF5gYLnmeTxwqaRoy/leGjzJ79NzgtenjgLb2da0R6iesLB6IlED1S2ehljX3NuNwVbf6XRsw
FOMozICibRnY1wZeKH1vjTpoq2043XMzXSbztB+6f4QATf8cDKqbOHR68/MvgX2RNXrtbwwB69VU
70fFh1aRAQJ3+jGOucZmVBD65OOoV8oMbv10FrYDxm743ll9JjupaacdHG46SF//NylLum1B7qKL
JydBt+yQRBeu1BR4rC0GjZTudI70Ojo7ZO372MyQbNRj7bzn45wrim4o4lUATMlmmzliv1p1uHQQ
n4xEFdQwAo6HSpd+/4woEjvFoOP57GobMot42t4+tlDjnLJoBD6nZn4t3LjOKJia+xSVKAQqJLwi
ePp5uxWXI+jvZrCuLeA+c/tmEvxboCcP1i2Cc1ndZ31DFBAZIjZlPrR/rdbKxWeKLZZtEy+08IDd
YT0gxpOOFv81DBvN1kVt2MgecyfqRaR3GzG64gtcb25eakJ+LMvzpsGB5JO7EQ2ONoTIM9kmwkRT
R5w9psVx1z/XWsFrRPcE3QGpe2FOMA2VsiT2g2tA52GqyTs8GDecS6j/FL5ZpYn+leUJ4t3ylHSO
z8eCCR5ADJGqW07MuyQEqvPFRZ7q0Ot9jXsAjJ2TEPTlg3e1SbJbny/Bhutvvq16lKB7t/lg1D44
VQhUvKJxXZQ5scCEI732kh+WV4ajtfhGq0ov6mj+oFdIzfqNYZv+iu3gD627HTmMMmAOkYk+5ZAh
eoJV3hHyC7AU+tz+A794tt4FgiETmV7Pdc8XNHXeB66U1jyIjxcPMH+SZ7/MVFSbRkWpm1LIoRjN
uJlA4EVYNQlc/VxW2m+5gSU820Qv+g0/0UO1/lckvenGC7ncW+ahUt+PPOyh61Q3oHuuuqyan85v
wXUdGrKayON/wrz383uzIVASavK4XVhtF2B4IAqV7y49VmR6kWhUNqO4yCZBgBl7dMlAsfxRzkpe
gkT4OtZJ+c/6YzXlT/njkxYN0AT38oqyWKk8VSo4KU17ye3GkccME2B0au8pecqPU1r8f8HuEsUA
Yh8rY3yVJpM9kwZR3TbF2efAiVOz15Uw29X5mbYNymR8pycPoXmrGJ+b7BIPCd9y28RRpGUns0Wj
7noR6iCaGBKEFN4PBAmp5JTC9as8FUCTLV1BFjrsodrZZRp8ldtZbcZ0HmaZMgHpDDh9hWkBHzal
++4/9rOsOynsobU1LobKY+oTFr/OrhruNvrnZ5Pq/iDCOa5I227tnPjaJwIkXC5717Yb7yfavAqg
h7WJ5JFuDW9lhSdEbfSoxEKDQaZE5Q516A1BckIkHxKTClAA4a9hftgOyK1sAvS2l2ngOtAcRNc6
/cKnRFvJ1gtbGyDMKRuV6T+uz/JmBZyVK5RYTxUz50lYNERccDAtfdL8d8a9kKCj3xbVWi2kS5r/
5V3SqreuOv+DKZ8TV2JkT/yvDM8VmfeCwBMhZR8X2X3Q9Jv/Sw6sJS2vREKgszd10fiFMIkziEcV
EIZPmLC3TYd6hOCrp7+XbVFx4MjM5O9KYDO/qBqIjhCd9PWcZHnOfU83BvANu32fuF48oMy2OMCO
1ZYYpl+WZV8do6m/E0vzd3+dsonhhz43UHkH2htinX0axyX5pNhJt7Bz504Bx8+cGf+D7ZgkOPhk
d0otxSyFbtASFDPAbjhSwyV4AqRRHZu/oK2+Dvx75F5jg2mTllM8ZFqaomay8XyR5ZmWCOOMvCmL
KK8PKP3hwPesf7zHUH0k5yOev5TmMXKpkiXXb0x/LvtG44E/+yIhd/Bqf+CBQOGQcamS5jt45Lj0
cTu////suGWCjPaShG2jUUPqR00AFS4TFKZCrgsMZcZ01lN5+menKZQwbet0sdWYEDqg4eaCq52S
5+lYn3I45cM/7cav/77vhuLTleimSZw+SIBEVHiFmpcOqcoW8LuQAEFZFv924TZH0WZiN68v7MnC
yEvb0wnWAqPVlyG4fmYRRavo3KLLBSyH6ur5q0kaeHai7Hqy4fIXJOsHRyXiLO5n2PutAO49X93L
ZvO+a1TopZMf6SKb3XhTveaIg+NupCjuMo7MdoAUpxfdiP4sLok7q3KPwypEJWZEQplfrkW6cUrY
IZ+j3/aKPsh472i4jMxikQ9eWmOPvzK1xoqWzIjAoE9iHjrxymMXbtl6Y/P5ydAT39GP7OXm5dez
xrU1PVduL74TjF4RROLjGV2pWKceO+8mVuGDEORdR0af5aqnzu7yl0LVuitndwPypMFU4f5xZ9lj
GUPJ/rZf8/srIpyP+AwiWUoujRcdFeqyTw9mSA+kO9c4vNgMEM/ZMiO64v/2ftN5uROIRQskguj9
cQHmV4UAwSmvVnKzWkBjisZxLdTu1iQCkM0yZvxChI4Gx9sHLlBqw2zGb6yy1KBrHI0KqZo1Muxx
yQDgGa5bIvHJw9fEe79RkncA+MaMSkynUnhHavv6QxSWZuX+k2cTMmEPsJKEag79mbOECL/E+vN2
iOR8hEmInVlWawbWZX/gsrxQm6Qk9kqRRSCU7RfI6+hoz7xhUP4FnvMaDoKFHSJLrIKL3MJ0PGHf
IWPYLV8Dcfu721X7TxKFUleB57HHHWvvdmjWNf1tg1xR2kcxZfX1P9KaLsK8ospr/O0eLXjcDvPZ
AaOXnlXmsCP6TvxV7SrRr46u/VKO0UnNgKfmiT48FuXXV/xHf8AfjcTqQqES7Rb+MG+X8WjJsUal
wme3XR4A/vhLL+ddZfkVXSR7MQCQVks6/70d1TPVrZ26jobw2MCE8r+0Q/Kp+3TX5CrxXTyYvIA8
TjqeonlGPPpaYm6XAI4MeEGtDzrQ5Zofdq5lQP3StRd4mWpE+uqtJUCquWUfIc2eANzzByllkAuJ
KDoLxexwO6v4B6Z7vr/vSfjPDQAr6a5Zq5Z6Nuhz5EEU1lk1JJzTCB9rJJkaClcDPC28aZ3hSjSK
7nlRaXPFACsOTHC0d9orIEcepwgrwWmungF6ENWtQorzkSaZLLcBeQhffBvtIe6mRb9+8Lt/nXjO
tfNSeW27AlEQEwBNmcPN9x9YGR/GSGf2o99OsmTyzqFg2K7OHvowEaO1G+9Z7cfU44+1hkXxmcWo
9AgadPDaGmKhN+ntXDHx7nT6NnR8o5fGHLhauLBURBkIfpKhpTgWVKX8bCnhk6rhQJcwG9eP5O9j
E+vTNY83yU8k37/BNkBrWCvt3MUBlEvAlZnVa7DVVMRbvqd6JPEb/ceWlm4wlnI681ZHVkOLnhDj
eOxBPJb5tlqi73LuQJzDOzbhpC7PEIrVUfgNM1NRZnX6ne2904LN3VamGH7YmYijE3reRwOFtJKw
2BibHukSTPWXricr2aSjkTUiWoVGcyoDg12RscKF4kw7/qxy285VKyP3LAhdUaZj68nYZVLQiwzI
65+iZVctMBIU+BAmhlDrj0GimEKFGrW9YIrQ90pUpG2gelNBk6iICLg/lmeGPiR8JSkV7X8dRsqO
BtnM/VUHU57IXs0b35hveetn/RddrcHzcUOe3kChhTAOpuopbjRWNvhfyQ3ja27VjXF94rADCEdg
rua9Apl4D1g9t5w5rfr9zas47Sc7+EhMukRdCX4WxrrWvKMPPTqwAbmwN7zKT43Yr7BqCs0W2l+k
RDdBK+l630AkCloRV8dMPJzGN47WTozpo4cJIoMjo2t3BlgWCeqZmZ5dxJSHG7cquCh6N84l35Ud
Udcx2D//97Eka+HjV2HoreoKW8KEPqn79Md51xPibzujA9tWpUKRwX5ONyp6IX/IRtu45od6qwAV
7yFRig6kN7vHzp3BKjo+sbA8s6t8KF/oiHXD1vH21lMgSz8Va+SAGkZuTBSciPmvpzhlJ5KLZLnG
JDv4PlnxsGfY6FAp2RZjtHHGCFOOQe1crFdUZ5Lq90FszA4m8nf9QKi6fq3r0/oVm3bsbRTkXWme
yz8KYgZ5aIerXVUI2utKe3Hy3UdDkqxzXMgW0czY2hNf33zCi89hpiKR5jHoH7g+wC6NeBe1ANAI
D1n8OvKv55EnIFhCDKV0xBWby2a/vTvktyGGJ4GfYZwK/U1/XG4hnYJzyRAHJAjwO1KKCGgu2WaD
yLNP+5Cfe7CAN2O48EsZSeIe0iuAndXMwG23kDb+Nlll8I172iSvdY28t19a1JfuFyLmztIEgtsW
vYCwEPqxhZPT851NLLKcPnvoh33CpQPk/grryZboVZSkDa03VStL+tgOZWxQA61KOikO03j1U3ge
JjAGZNu58E9xTj4nk7db+IG7PW/lAPHZRXocvbt02s3Q/9MAu5uCip03zuzSmqi9y61cqLM6BAwo
QFRc1QVTqj0tKS9kiFLQXzeOW5DX73SWxliRFldZ2bM876cV9vxcf0UVMVSZEXsX5BuhTHtb1r2/
RvF+raRLeCJTlbGdKviUyRiXlOS5RDi07iWsxEa/klQUMjoSVgYniSPGHS5n5j7PK0zSnDw90vaS
w+DeEzO1D9roEqS/KVmTyg3jIlXWdPBODC2WkvOsOJ+yAWL2lLmHCvuZnkUsMvY536/6E+Qqo3LQ
RS5v+W20xGhcwuT+cCqFyuMosUAHKMdDu2DnITUoGphKdjsmjvosWtj9fdrIAY92QrfCZJaidZih
Acz+apNWfZSTVIwJ8RcjGxaeILvrTXxnL4he2RMnRJMK3XHaDnQOgo/sNog8WOiDs0MIoXOVozLS
99O6rK77+/B63xlJmVPeNwsqAePWAv9IFgJF8MZDy6qh4MAfrPD6VwgEFnCyuboqk/Y2o6l9E+P9
UX7KPZdhAWoeWpl/lZvLG8U8ZfRLgy+DlNglQaxebi3+tWeKx9jZM1hDCHLEFoQ2xyGOtiVY/VH+
zspAe1+SVz2ohaqpjKe+v7EyDqCD8uSKF4mWw2ZQ0S2VXZoH5iiTxWubl8+clABb5PvghgpXT+IF
G6D0xjaMGLCq6VXv09ajPo+zAvaRCNZL0VX2wLEQpVgyvV38hWdpmwmFDKCp1sQH8/QA6rKOR6B2
IPQQlTZTtksY92nXPsXc5NTCvxqx5v3WLYywN2qm/yHh34nzl3oo8yiCRvV7ZqwslFmupRuZJijl
5NnVAUar/ZLbdiCo9/lwSL+G3yVpIwF/VuESCLbnhclC0JsonBPF5jNH9NrHk/DFauKByeqSCH4i
79DJCTsovkoDV9AnPgcv+vKu2ZH28DC3cRXY1Zgumx3QMfRO2IqMrxQsxDOJpNm6vLKNJbefmrPe
fOS9MG8Stn60NCMHGj/diJl8lvfa/e8dz4njQ+DDxlwapTdX7vsh/mC6vXbHKzB+lidyeoEAlnfA
VX15yW79cJtTs5peAcjEjOhiEahwa/mbosHhqJg8UphPG3zeuAEqEfiRqZMXB4jRo5MYagZwsg2A
+W6mTwhxTqRHsIZ+PBPmix1vWgvqxyLHyOBK8O7UEcm+ZBeoJXKi5R6KNTnQOmW42pqPzebxIRfc
3DRXuSxe5Hr5nyMVChc0VH7WYgpzXEIx0B6WSPQcYblnvw4x4nxlBEOM/jsy8+AGousMdmK4bd6Y
qcJhPxzOo2KSyxMtvFSZQBJSBLcegb7Xv+3yrgjyJ+77Mv4V67rwGpz804gONNMOInh1Ewc6mTu8
JTr9b6h15WSH9PDTus3g5uqCDd9hCeo1dc3vxH55EOALJTbHW/7oIZNk0pJcFJC5ejOncYcgQgNa
Qe79CEoIzKrjbzItuim6Wpsu0eF6R7vTaqdRBTawcQxH/1JX4hZ3dAt8MpSKVAKiFFpdKGOLWVyY
e2koWe8Xo2lfq077EpmBVliFB5d9fALS1z23Zk6w/trw7S2YgvrkTfP+Okl5Jgu/tU+dzyuQsvt1
or75zhkmkFXUCKq21n3/ssfp34WWtRNTS/NE0TIFrBzsMuuMerzSRtMnQV9/303lD/8Q+iZ+xMwW
+uLMTzVFqm6sGf1/Z6Nb+h/Y8aII/mmvY19wWiSgzlww4palzLylNrmA7Ah+wxmAk92FtI2AKmpK
r2jQSN9aqod3bDegKEDpyTMuj9hoMAS+QQOvsf9JF7cbfSqUsQ5LBIo3MGFtOroIoI5Tj1gkwu3T
N72Go0eGvjGAtRxAjegcZ8rfwFDuBFzdnolzYLcDMpIrEq9ZJTS226297SuS1iWQAk7nv9Cj1y/e
GxeDjoeS3RJTuqr7aLahN7F6FBd1ob/J/Q2tLEeusnsp8NY6FqpuFGI7weFMWrVbavs7SvZlaPV0
POied1HeyW0t+kJ7rXjcR2+wNbXVKc7U2qvroLoaaub19tF3k+sSKmN5ujkVrsnVDkdUqSo1pWWN
7TsfVC2j5KR7qVjgDc03HG3OcEiHeIL3xbesGvRYEC1Lhe4oHY6+Buo35oh9fQVEXvCbeasWl5tk
zyCdV/L6BCclW+yb0ZT9b3VRW7bhi3XDiZm4FnXUJZ01aC/LOUu3cjroKbV5L0e+QpLZWcxx9vTd
TSgnd0vFwwGz62hcd7+Ondy6UndjT3lFb7Ha8MUt8xm+bvaS8BfeekIIiF6Rnbb/m6ILqyg/3SY+
3vH2GQQBmSPGBLmK4vL6uU1Y7brP/Ju9cCtoSLgY8zD1ZphPWiFPf4tNnwGmP4qWB4eZJYMW2ODO
6sVqSxrO6LLNNI0BTp+LT1WF+Tq42cz6cqFmaDALYUuuWLuzrXY1j0jq99UjLHLUAhwEW+A9zqcv
D2739ikPZGW8c9b4DVVJ13JWDmty+hS+y8SZbgDisNOSSDdwQiD+mKc/mUDVHnvqzQMfCqalbm4S
KQJft0wgTMzb1ZF8HRh214PWLjEhgaPm/5hHC7ddLamnf5rNAhvU7G9JmL2POLW9CTJGW8fzFWP5
68ob/4k+gP8YgNaUYFRqAe4KyLNPz3TdeU/vQNMvI3XcW9SgjO24KZaClzTYXxRF0MLoe2zyIK+P
8x4K0yOwRV2RvZDmPqRSECLf6JdpYU+/Wh+ucORs+KGkCCniB8yrULxvPEhpM6r4qKQdxgBiuO1B
gidvtCoUy9MdrSAlK2NYKi/tQ1ZmEE7o491mDslLiCNrUg2k7kG6Ea5FmBNnRCfMSbFgKOFFR9BI
iqgihiYBgDa5tfTjutV+NccJVDEmkYQZa7QWdUevB2LyY5e2C3abxvmX2Zb5Yps3wYEmmzssLFHL
MwACzt8kQHfV4nNR8S9a1/fBu4n4O1Qu7ZO/7Ln7x31xT3nRgg99G5xW6a4jVG58lj4qsDIgQhoz
mAmo1kaqgU6jr1Mdc4JdSLyQdCLe/EkJQnDGT1SzfLEqYnJsISSo2zggqKQRkYLXAIwbCufeMGmW
g9Utf1xVlCf+HPfJH/9norTefeAtIcc2oq3TVWfmT3PftJQlcgZ5csy9RdbjDOCiF0n4VRuTM/dQ
FPAo4kXrlQymPsaCPATBTnNRGMIxeK8v5FjF8etpiZcvbPT2c4nQe18xjypuLw9R6xVMNA2a1ROs
v9pIBO9wTVKrGt8vrqDXp9Hwe5P5+c3PMfAegcIHcXLr/atRQXziTsuwEcpwbrReOiDnFGvgou0U
ekPAGlh/fa0XNpqJpdKWhVNzVO7FIS0x0gJuOmVDzq85X2iNV0wdewD2H8CpX/ZBNjbNJi9yZUs2
rRwc/4vA8+XCzBzdOvvVw3Sr8jMdfbaCJHJikj6MOzm618vaSoW19nDSxdjrKZq5ixEaU0yiqjmp
CH6+uMOttTwH3lkb+bW9xx2r21hQlSJgKs7epcCayF+f25dLqxBtC9heYBFEkdST9fSmIYmq92x6
0ur/aL5nQ5b1ZJ7CpcYTRrsMPZ6JzsLVlBXr8vuLskl+H2ASGfmgEw9C2p8zDGrm3BVEFPyiei04
bX2z5M1XB/SbDQSH9cRQJNrrTs+4CvMtLDKeSr4eGD7NicggTR93LNvBMUOoEWQGhNHb6WvSlbcX
UlJ8+RfvxzhucRzLQ1gPQKuomNN4iJa3Ok8Rv3rdm7TAcXHRBJMTVwJImM4vuISm4yVkln3zRy6N
24r/rQy5UVvoiWO785o/1aGbgwSez5RQ+p86mTD2NWM1d6Uh6B8q12V6AMiL3aWNQgn/PZs2gCO+
dKaFQAJ59QEzFo/AqPY9FqWHWUVDdytZMUHfS1uH8jiKd1MedswsSikUj9jWmvKMQRLuBDdjIJHl
+Umuo0iiOz5xxhafnaoIkhCF7Pk0/xGOeBjAIKrUXEkPG22ej6Z8DvQEF607mWAJ7ONCgkR3Ehws
geRU61ewCn7flAAE5LU68NpsGrHSaLIi8dbDXY+xHY8NKmWKjE+ZLBtr5Jiz+lGd1k2DKa+w/lRn
RcJXJ1ZLrrF5G+SMhjiqt4oLddXZjJyhSqWEx2y2IyHRPKeQrl2jrh2rC9cYZJOdnDAUY91Oq6K9
07Gh9TCLVgjHryLgxzCAUMsPWiyiprSpmf9yxWNF6lrTMWrP/GHq/d7VcWqHCLUt2hzupaleaOEH
RaML/IU1Prn9bSa2+0NQAkKMPuaI8JCf4hnduB3rz2hJqQSqjy7E+113i6AiQh9A161ev9YL/3Bc
b7zIaEFRSa/VwdsgfzwHVbTXqVunZkP6Mq40INS7sc4uvD0Vo+pwLhdhYl8vJKH+YiRqQz6DtuSF
qdvSl1ZauMb/9SV+F85tHTzUZIYBZdmJelxUjLI7UFptNR8N16oi4RekRaLqY1eNlNLytmh7H8Ue
6H0550bQ8zdqPVZT1X9Bscnq9JMWX+SjYHIbCoOK9Gg3mhV4G6qyEBlqIkRw0IIxIxy+ZZ6C/81C
3BVp57Kydy+Fn7Li3/yjKebQPThE2yycO1422zK8F+E+CESJYXTl1JAgAkh3PR3dUYZuH7PMolZb
oRnRHkudT2t7QBAEdl8dRmQb2U4OqSHIw87d54lqZAF/uhWdyoV4Fj+P8RqwvzMacRi66aaHldMd
rCmkU3YdoVLpb1bwTrlZKmQkqtIMULmltGhEoFWf0uCZGHUrlNwaIWWV33fOe+TREYmTKWPHhnPN
/RURFdFQwxfVno99+Z5uLCNEyEmoAolK0GxkEUTbT4FkekWRVHQraaqXO4/NxgFsrT8qlWM8odJf
MuDsJtrhX5E4ww5mv0jIeTrqXfBnsviXiRBWsVLljcVLX8Jq57OpXHC3qhGfUHoFiVoWGLr42m3x
IBqNhr8u2M/LqlnNzJB+PiTvREW2ruGQ6LkRBvnCYwD4QmxTyxRVAnIVvHfYyleyAQFRjuelKiAL
r2oZqeaoAn1rGA3VXsKTeaxXAUp9G28Ul664j0+Mpaewwc9TiVx1y9qu7WI+hceWFBOe1ubXiEsq
2/YvWvqOjK4Bp/CRcIPk2AcRTNYsdlYti31HQfHKjNlVVco92cWjLWaIv3ZQhzOFL8ToloaS6D+1
9FtU+3aulUs+hZrYCuBdbopcXsdKBlUi6a+i3TjNymfp2l2s3NODttxGWwGM9rCVtC72Lxlgtk56
zs5fgNmC9XWq3TuA664Twt5W28Kgk7U6zO/5I5UbqEogGr76H9aWiQumefCP7p1tcSmuYKuvQlSl
a1fbPSrkM1YTw4f2bt2NSJZ/Zog9TtogjqexbyAZZIYj0n5o7b4xQy6yyYhqlCpI9HKdmVi81nPS
yXAgIxKjsg1o2b7F/cfvhgNRfjBlD/3fVrh2OUjM+TIGsc/MpJXQBDplV+GhT9hhCJD0yovVJs8l
BmdmoRKCMOUG0RQCyKUi882I5roJIhf9bt6ugiUNW7619TkXRqbuFwjI7O2fKDrvO3hgVAeS2Ofq
pFK4uxWdT0qWl/MnwBOB1tE4RY5ZH99QcJAF4liDGbR7JGUjGJtX7OIjQuY11g54WmDJFakqska9
zKH1F2j4ivipLCSAOG4yLKS8q5exO0vbc2AhWk0IYmLg9Y7dLyuOzHKHG1BhMGF9MU+DCzcrydgV
FZvgXagoCQYLPq9cF0gX7PGE6wrGcFLxgRP1CJbFjOpYU/1fVF2k99c2awTBgHmwVFf+2zETDLRQ
k/gd1qDhQRPyA+ot40uRlnk1jF3GYFfHDQHXHWZW0+zAS3qel5d6w2ZAQLjIo/0P4/osIngglL27
gTI8XpgSaaMjfZzGtv7jfNiq6zhENRy5AVL+1KJzTJ4X/J4blYu5raetlr+IwR1T3mWszgj+qEVU
ILjDVJZnwvqZFQoulfZ4pxTZU2eZmd4qpb8KOZYQyuy6inD0qh8AcqqD0/tRbuqVROOKodDZOztA
gD3tuEQmdxafPCDCfYXxv5QSImEVzbTTPENhHTsr/t178/2NBv8caw9h2+fgzEs8jKWqQu1V3pSX
tq3SPDFd87fuyFYXKe5dlt2MmEnoys9IfYOitFDboUSE2c8n7Hto9xmzbpaPV6F46B5dWGeS4PwT
2m/xa6RmdghtAcBKNE0X37cnIyrcrTkN3hB2luecvKyy9LfVdi5hDda2o3RHDS8cBImtwtuKFO0v
BaI0HqmaJTAySJ9dM0GN5S7jeNdo500YO3uRwMz2swIctOTtVXDwZW1ckLcdJUcefNtb2C37RwNE
3PFI5eQqQQ9A4z6RELyP8d9PlC+I/uUqj5w9SNbA5U/yZHSsdji4bSsWL5Lsxe8aXLebYclfqNto
jHjIcP3ODfZRKz9PAdy1mgT18uUUEWqCVyfhzRG+7k0zyL5jpUEAADGGo1oQE+ts/+pF9CRsWX6O
VBoN2qvHQ0tAcPJporu98C5qefxm4fSymuFCJqa/Ine9fLqoeXuTqwLouNo8UtQEbupQ4ClMLh0b
wNpl4apuLDLar/XKFlHI1fWn1QZvGSVzBvDIFyYf01oFacONVl9tVne8QGtPCnjBa7dA5hdXVz4h
DyTDW0GF0YE4KIpzp3eOGC4Q7KLeDcxWXSYq49kiFjXUDDly+LXSL9lNJFOYjg1bY+UHmp/UeFxr
tSLdciGy6AnIP6YxBUgBQ5ny7rClDDARxrpgSYmIj9yuZHavNTm4gg7thtNcxNpArt3myf1Ape8Z
rB7jlu34PHp3EVs+IuCtRYVRTbR6/kcf19j1AgLM9C/CvdXdcrFwEOq+P9zd0ctU4IDogEcoXmaN
zj52gcD1UM+05eOw74jcrdm/4ZSCiGilt02/v70toQdCtZ4MbE5CRWhXpyZkd6ntp48M4kP1Iq5E
A3WcYcVjX+qaPWuVo8J53o4Q/DQKfGn878dt+bfsb6bVeWZyk26nqtXj2b+qq5svA957ljKXbzxi
cTI2SPewhi6yaQKx65kc538ePJDk5FFXaxydTsyqggVRFxnWwJVRlgOEbSQQ98m1TsTuFoGdhz7s
xlYfL/ltBzLnH9QACQjuE6Y27TUbAf+csqdlEoDVzkPjYzyc9eaUwZcluIOwlmgslu2WvE2IK9vN
Vl50CWSOfG0kbHL1mA6IzMub1QU9q1yQAgt5J7qfJVtx35kURMI7XvxN/hSmCJy7GaR6JSVaCVvD
Y2HVCdmbSdhcakvainy/b1qnxb2r+8j+o5/0SRAXYbYKkDF4ZoDheVw+2zK5IHLjyV1cqS12KFv/
uYb61ovbdUZ7gzxlyITvDXtvBjqRznWZtPP9EubXZxnV0Hk0YVCCk9N8xfGVId/In2X0xSru+gHE
ChpgFfnr3PeyNLD74rbfzJMGVuxK00480iWwt7lSVC6HnkFhuPR01Syd5xCzzZAhV8TfYfW4Ua/7
UdGOhalZbVnyCNcR+lvNLYv92vzK4T88+qZ2wr3asoCl8iup8R48xXGx5WNM+juOTGMgK0IMKfV7
kW3pLwq/cpydHriUaGubYGrQIHbpzx6PmGzPIwvBkmpStiwMBARm/WAalY9sfO/L1BLSLORA5Lm5
ODmK6MA/QySH5hsVyUzzA03K7RupCOvepXAS/3PMNCauQia1W161QyhGMMwp5vWfmWWpzRIisg9z
PRwLYYjgkyqWjfC5GoSPGQJ7fTe6s+3P2Tw6qfpsveKQwLoXS83p0e0QiuSN4vSUdMSgZRWlSKfA
K3jEG6FhDu8lIXzhzu6IRcWFu5+qqgrwyirvr8zW9IqAyCXKL20J50BVkFW0Az37yAanNAToPJI3
3SKTqBk++IwJaJ404cGcCmKdSrhDklkKfmeWNmN7lZRrJxHtRu63Ki6iwIXFA6ylQffvG9jZWGrl
cpyDzRNIctiImgKru2veldJ4ShqpGRl3Q4QrS3kdFZWpvmx4kEpi7trmakKdfiClMUvCJA3ZfuyI
niUmg+hL1afsl2Xw44zgz/f71rN0shvYWgtS75nGyA1Hv+/n3otrljrx6C8BP8syX7tVkOimKDCL
tE84p4veIHZ2J2WDY1xS+z9GoSD5JSFuWFnf+d8ol7dK8YaAmVIZEMPDGXKLrzF8lkLMWn39UVsZ
H85vn2jMcdKeH5op+pEmDbUHoDQ14sm4ux0v/66y8mrIdtjuPzaF2WU+b10qL9e2eS5VH6SB3E74
CxnTJciWczpc1cR7sM6FQzw387GSeze32cEEq2mebgzE6o63LPGABYErd05E/s98amrdUxSzutB2
5ON52GONt4XT0/EghsqrsdqIjb6CnuQPDyO3RCVUEk8KO3QOmIjOvB0uUAri8ZD7aqkrbhk6VgYl
Rlyxh6Qvu5AziWRaOf1Hoa9TqpvWzHIfJhDOVk70HpwWPnebvewDj7b9DaRZFJ0rBTPPy/DSYyOO
iOYBKZiVR9UBa7LeCNFUW3r9cvCyz0leq0lVVEXgUNj/jr6U0k1No0Cz7lIEPc50mBwzRz3lXBss
Vb6pCzAhy4l96ax5C3rGWbTlyDKkXkv/NDhD4bqAUcd8z5RzhOZcN0MTngVUyOfIRolW8moMtZKR
YnpJ5RTDODNvuDb9hHlysonyLjMhUR8Qcru749FhqXoJQw0Qej2l6oMEM2hFg5xgwpAsMYPMswcG
mpd84ETyYtZ0Wsczl6NTJ3VjnK22+jzPYP32motg+rxS8ueCc5tSpYEyJKj3ndP/FsJiY/UYQ0Eo
invDwsdbzMbPQfd1pAM2wfGF9HIsSq8uvGgvEHlj7Z/LAXGg77e4J75sa7tj8hcTx1BGdGH+390W
lBujjN5OqEsUF5ldGvnegqd0i5tGCWWE4vl1nQV8arF6rSPxHrThtD276eilcwBNnKJ5MMTdzqIt
/yGjvIkXqv5zn34WYKTrBA2Thh25a1dDUHXSr9O0FCUL/77IcwRepRzWmjzDVFnvukO+NG244Sed
37JMKPKxWUxH1SYKrW/gRAFrXVtWWBmlrqXtJHCaAVBR0HFJTvBZjcs7tvmZ9ziDl4XNfz+GOLgz
ikQvmoMRKDecnbZJtnj/+D0KPTeAakELkT/WJZ5ymHKPl5LBxUS/GJtJ/016vlw5OQZsmJ5cxDSR
fFpUVO4Q1Jd9KhzOQ/nRyYg8xErG6vWRKAPgCf0Oi7UnxQzdH+zdx38mnAExstGGcmW5dtHxH1AZ
f1lPZuTF3J6b5ichAopB/0lNYO1l8rULAEsIUTyuQar40Vu3Pa8jFVAYvVLI0ew+R9v2du2QAJ2M
TtPQZY8omIlTD77GrU8qgM26bI3rTXhV6OZl4QEKLYZeR1usFZ6pZU9Kw5VxM9EqV4+XMPMnwYOd
Yyl5+w4ZUh8w0Glw8vZG73waxIDzdaloe9gVi2uI7csswdUHgMQGRflZqmZUjqvUwcIeO3nvpb/O
6ibfAiBaO0t1Qmes8DK+3Gri+CwzcVssPNj2RnZgaqb1ydLllS2zG+6mLCh9K+sfVJGiGK3QXKGU
AewrFdGPuxUQ4nrbcVJHKCjGlMIZo0HAPGGD97CQHnTn4YlaxZQJfz4f8+AxZtHb0un4DLZRzo62
5kj1Y1nAsJezE3C5+rrekzRmVwWUI9oQQjo2vCZ0Nko7aIfp/yOoyYwZQeMR8WMVfPeornu/HdKD
LPz90wLzH4+wNYGHNgNN9dBfl8poolKEDEHHSdrWvb8FdrOEj4aa9VepM2+sIraP1fko3OdUSX8E
+K+Q9qnvjR52M8CpQVfTY+3KDvqpvwUz5llN9azYi5XOkCHOwgaQjVUiRN+qHlYHFLf9LinygQea
bouqsq48xh7jHMjgZevzZ+7R8fGBE79Oq6YJcRBB28lWZStv7OGjLIx1Qsn5rWODqH1Rbc2jgJTH
OAUVV/MvXJgQGHQvhL376OOc6xzTH5Pfw2TMhz+zYf4R9aXj3EocPdZ3B5LE0WyhwQukE3HmciHe
Pu+QxvUCvOyzVZsVaDb61acsTnNZRlYziLRJHHk0yRlaS2rES9GdVl5kh0FAWLeWwLSAzI33g0qh
yJWbDwF02u8AEx38D7yQw49wU5LOg613LGmD1SonCqPiHGmlvm+DY+5r5qSmRM3jT2SgoNWbdTji
xLqqmtLHJVxKaYhHZK7xKVP9SKQhUlQF3Bfx7sS7g8axcFB1LXLCpZAvyPAWchLf8E++K/5pSpoH
7fW+QaTTTI+QwxPyYnpLOi1v8kHIsgxvCfTkiJ7pvFFweqtrYnbTtyg4RaFIobCqmIdX0rf8viUg
CjYLM8CUuIM71eYAcOFYUCEwM159glrdLM183c2f2bpRYxPfjM5Xa3R1JFjo+3F+2mUJ/jI6bO2a
0u9ynY75bpaxjdytYKhEvRByPnKtIPT1FSfjcthUyPTioVPRRcMU3Z950VuezoukS+Z4Tb+q7xFm
Q19yh/K7Kg8A29am7AwRO0skdO6U+aD3NS/CPgwFum3+3SEdK1Ch0FPVY3nhVWs9fzY71XobsNmX
+uch54L3F1UaRCQxwk3MWUscqatQEriA97dod88CmI3POv/orEc3lP2Ay3uzPUDYCPpV/vHazUAp
M+qStTvmWrKmqGnKAsedufCCQ8eRzNdzQ4DUHg/Q8a2UcMgm9a/Nks2HwnGQa6rpBDR3F6Cgo78s
r4Ni3zANDapD9f5i79LhasPf5ROJRfLsSnrJD/6zLg961FsBp/X8L7CtyM0zjOHZ+e1LhXwGrMpo
l90A3A1I3nU/RQKC0VBbIWGMkNzQ8tEJKd1MISkR3bM+qZjm+gFufa8FDAI1KMtxCi53EuBLr4Pl
U99p/ajWTlU3GbE2eqvUYzCcQGmvRC901zLowNJowef/jUrOoWzHI7HjC8cgedavmJY72uS+yARP
8cm0ePeXhdeHk2bmV6ez28oWb0Y53LEW7bBpHY22Fmkr8BwniimwKGsFRoz5/NeKXpSIbJJODgnX
cnDjSjb2EMrG7TRn6h5+1DaCPMSluzOPcOfw1VDmuGfx9Dixw1JINrVw0uGYhpP4X2F0vrxlEE4v
SNtAaT6oWD6cgHmJWbaFTX2gRBWBEpdSLAlJQcig7RgRWIhNTL3jwYvtrlFQ1/F440Gw8ULohgcX
U8Sn7vQFd57RHYZ2TKS3bK5dcAfKdltz/bVDYB1ZUixt9wv+FtlI08aBa2wom2SyoJzVIxwzU0Z2
yeAW4bGN7znK2DXuQqunrz98xp3aq7tLhTejh+5XwX1BCCgiQHEsvKg5nznI7i1odaeeBk2y/oOC
FRL3JxWG5TRVrNbLb63tZ+SNZqbvxlxjE+JeM9f+USMrB667CkqHzEKc1AaW1UzWorKeqqF5oLWB
/xcDp7jIJbH5iwzHDFqeWMwLEUlb5vbcFnAa4b5FLciqJuFc63kFl4ZpU16/98FA2B1v7Y9toRE+
QHf9XTZhPQDT9K2eqXzZlkSKfqDGr25TU3PXJ/BoRCVt4/E8wFHEx2VsD+SZS90uJKDjrE2P9yDH
GQP4C6qY6tQ2gHv0lB7bGF9HcraOwf9RxqYzqGqKQYjrDcKc+FM2rLbsl8lGswTL6uL6WbGXwhXn
EQ5YXp7kP+jzisFj64y5CxG2mTuCtlgusZ6v6YydMc4DHFwB6EXavkBisHs3bwCNQlTpBStDgOMq
/LP0tKcYJVA9lYDDcs67DWH+fmOOtMNa+u9ZmGM4uYx5SjfWgj9eWVNlmA931cIj+t0/+GIvIgvj
1tqH9TZly1dgY55xUSNwQXdDcXITW6UevfRDJwz4v6FEdDeGYl3AFS8cxgxdsBKcRXS5Lsq5fT8W
m4GySD6W+j6x3Kwu7/VZ6Mf6xrxzejluZ2eEOmoYCL0OQgs9J2y/ZKhKF84T/0UspXTgfhJvSKVm
00O42sHxfE3rw7wBN4FLN7MzogFhu+v+hjDxMUB1ZKFGU4/AdYz0majzS9gf+WbcRiKn8KrYoe+W
5D45ta6TwjZVKv3m4pHogdqhuYX4Vbd+K2G6lGMSVD+xn9p4AJyEjDhYn+Td6E8s0IjxieJm4HR+
UJ9LZU7wNvasCUBjW2cn+vIznHPQFvhO63HkYRKpdKlS9tGQaB81CsbVNu0IXmQL+uE0vnb66UXx
7MiVjzdYG5IQfOYjOrpc8kyOiLXyHc0al11VJd27p4ZVS6HigmoE4UoLAjqWgssMdhfCpoEKKkfM
HWFJYcBYZe3po+/vFBleEeuwdWbfhg05Pyjjz6TIvzE38WXt8sOCtk0WpiCxOs9KdKv4hSnI4sXA
KolwyTIBlg8nDNULBydxmtDixg9R96NEkzBRCYAKhEoC19w8rBh3MhkjmJr2yi3qPhjqQEWkjMVY
1FXC1nlkj6qifzGyUckHckWNXt+jhj9MppbZ2FeRIdxpRjJ7Wv+4CvDNwM5J7kwEHHjoRU7yJx8b
/auBcd5UrclbWk4nxQKJxfISz2l9OjRPsC1RNwqTOiirI364VP6sbU6NJGTR7vrZFJiz+nIhi8CE
7htC6EE1u35HPW6etsSkHrq8I/0BlT47ymYyYZn3s3OxtA9Ico7Hci5mIMA0kvwFOQMWkwWPw7cH
A+OXmzKE7PtFT7q+cPNdOW8Hgx5pP5HwuUyBqEMkOWaLEeKEt2LaXJi9WDT8VfUhIb61xzbO4qE3
qd4BXp2LgvwiO2+CgjROc3oWu36TkgjVirKJVhDOxhUcvsHXZYvP/GrW1rbiJj499BQ/xPxNh7Tt
pesQ3R1XUlc5t1Fcw8N5rDzYcXzbiilCp+mWo3RQLoK7cEQaZPeRjCfLnwZBBSGN1zb3L2UZSQ2h
KMvTFP0aSHSqN7ophK5x9bQpjFYOt+W2uJUv/4bYpdOY7zRPdMBkynE1JEetuRjvrhqx1zScao9/
SB0XpdN2tF5LncxLxenPibCEFb52UUtkaRlira3ZLf4S+y4AovLnQz0HJFqpdpgePwxNF0HLJDtT
QsQkjucPaYi1MU3Y1SWP+AfLBJUHhY0CQmi4huI6ZMca4a5e0jAubkUGvEkOh0rrLaaEe76W9wJG
GcrNvZY1XsNRm5GmxaiBkcdlrvemgasmmMIVEb9sAsp7yog5xqj1C3h2uFAFBTa0VfVq7Zc7o6u3
sE+l72ze0Fft0w2J0WsVv5kdu2sVN+2DASm/TkhuJrBghNhUa9FveknazsvTz+Uju4DDSXkKsl7O
pxyTiUdl0BhaHTmNqQqqn7hvIm0Aw+870ljsYYayNKwGBWGaBgARc+pXzYgmMZ+oqYPENHXDHdq3
A0vILgI/mWd007ru7EiH1CyN/HZjYk0hk2fYQnc/H5P4kAin8BJ0grov/fdHGXoftiOkmRQHMsFs
HHBdP3kYWLAyk5denq+zAM/USMjOEfBAK087Ua+1BmbypmajRXEU0XsUfhvZx31YRNu973E2tO+V
4g8Hz9jIezC7cAHC0QoGxKydI4SZrQeMhbFNJj7qxmtYqiIuY9QDMylie/i5Smjcfn4vYYDbfkpn
aUu4UsdAgD1nRANzs2XhRbviqHtuMIkPxK7nzb4xne7djSh+hDu4SBElRdFBcFny/KUKmM0GC0PU
3HYXB/0W0vOoCgiJKvGxSqZfYPD2LXzk9LG7tPVIlqtKnYQp/F3fviijY3OcoNvGyoJ3WsBS6O04
SJb58uN7a8jc1bsoLHPycmev99CqgceVq9mNImSNttXVDMuGTF1wZjg/Igc4alXquN1zB1Pt/lXg
bPb5fBq+hGPGLcTNghG5PdnCUSSFBjIJcSb0VG7BySTP+2s5Ln87l18m75HNSOVzjwPP92toOh2t
9Ei94/f8CbHl8DtBBhJbwIF+vqtXMGISExE7BvJoE+t4XLltlHGnj8yCkgKoB0i/vKF1H3SDq8wF
BVEVc2R+JQuQkxugavYTqoZLc4iqybMemn3AzSUPXwsYa8WoR7RcJBT81iCZuJ/PrCbGXR8xpkF+
TseaUPKFgFLS7vWbHx6UM4dnuodQ3zU9KffPPxKDADULMGdpdnDSv8J0SQjClqEp2E3MUMUoVpRq
p9nJzFrwgbwO0v8biZNL8jiroI+ZzwVGmrv9GIfcSLImyhIs0Ayp1vQBnjPPJ2OogGXbE0/yJ+sB
yEw5ZkCvp1cqiQKIGlgRKPs1xpah7UFKmUrW0S4q6PW27JxgDIVQ2DHlNRuEkbgLvHhQEGdBuPNR
7FAEg1vjB3bi0o2fJTweCfWE8EWVBzRVbm0my4zlnIsIrsBM8QdLiF4odGpRunEKXXQ6NUCVJTmS
0szXuaTayvZ9GieoT8JvzFA9aTc6pHEyQ5M/twHyBUdU576GUffx8E7JN8USh/l4HRHZpjPA2WGQ
NLl7xbBv7kh7PnkhMTQ5ly9lc+jHDZjLqe+12u+wzOx2gXGB7+FfsmxyNHUgNid0XwjZ/GMvxaDU
dCL8oC4ZNrRN7+RRVKIyVmqyXfUDrOgL5OACz9CqLJP0BxYTNBLP0twYvQHHtqeoA7SG7xkdZI2I
8CafrJwg6JNqxjzq/BQXJ84U7JgcvVFq4wT9+j5bWjSi/CLt9CV7HtJsWouMB83YVJVS207YMmwY
7GsN4hhSJaIORSd10FLdCPnMSGW8D8AOnjDUTIVecBhN57T3KqSOh02LsYQafM8vy2x+sXNF55Bz
ozFqZCsSkK+hzZYZrpOkM6D/wa7W0OTR+Kboh/ynBNnvu3Znoq4BT4OVMChMBioxkfpK2R1l8GRO
TLs5cN+Kl2VFbYBuULSNI/PA4y4Q/wDAAM5ysQ3R3kHsu+9EPkBOKjsFosIHmmVIo9ympM5srd0j
PzJJeJ3bRbHsPNu59rH94ictqiiyluiePCdrvBEDgHEMyTOR1zBfE31lPDdvaQd9DwUtjV/dacYm
EjhLxTRFDHZ2WFRopF8ymWs5cH++RpNOkQnZoOhJzStDhe2/w8y6GkoDeQqnycZPxs1qhrwi+cms
q3pwUMZ8IypV5CZ6GSUTo0ufsnmzq5PBnlUyG3rokBq6cRiwNaGcCzwBC8LDBAhxPpieO0wXXtWE
k0LbFxfSgdAiC5m4njoqcJlTEXBp99JH/TZFtwc61zTgU+YRh4X2D+mrWUNHyZybQ3Qn4FjfDDCC
icmGAdo44XZjAp3VtpM5HG7z1qM8uZCRZXHaHlIykr1EEKWriR30jDm7E4/xrKUDLcnLHrZopmaU
Z865OBcYcVznB75o4gelpWS87iybizEh14HDM273DLsGLOpLfbDOGGUS99w2jT819409Blw1i2+T
VOMKPfa+3uvBJI3iZKzujZbGawQn0eDKY6vmCLkimT7I8i0sLRk05I4/AUNIYH58ASWNApBlunFf
M7IEgAKOi3j/bm2K+lzJ6cjtmzyI0ZbLYWtgZq5feP/WTToAwFp4Szu4T5jET2itX4cPpNAOF9z/
9D1GmRvu+yNrbTmMrnsiqc19O2zmgtfeK6t5YTrxVg5xkxx5omFkjjbyqP9Bo5J+JeEYCpikX8Xe
OJT/Td5xr5l5mcFBxbo90VdG4A34yhcHT5JFn0H8Vk5Kdo18YKgGBugtR/fFnvHOpodAQFkVBiiz
3yd9fat9QA3tj+ZyPQv9E+BaRwaheHR9ZxwBBmQ89PNRZo9kr83XfKCakioQRQzAUjMZNv6uZyav
/iDohWksmuPstUUfGoTrJoWqv+3z1vqBHfcXr2WQg8BSxVSH2H2mTA1vGyeRglNcZugu9dWy2uek
Z3nknawNh10QDBiUzy3ujU3775zmdxmJE5DJ2EuDJcRVS89r4v9W+JwIyE45XAqnPE+7Hhq2lhUF
1JV1micUso1hPhIA/eP9hu1gh2n9MuSYB/VjGEj44w7ueSv8JYj02/TUpAWcM28NU3MV0F3uubol
pTti14owIMOOylY2fQPAiWagdR/0ZukaCJXWBBKUiHi6RPkiGcMpfKTLtJnVg6jFGBHVOeOWp8D8
Henfmo5ytmbiKbObkztD5bszxliR5hEVwL5YQk079MWtjU1s9SuMOqNH1hGp9SkAxmkzKZJDVGBI
CJP9qt7ZaFpA1n9ASQJKN+2PtMW5kHwhnh6RwJV66ZveqRxCebwmT1SZu2tVX0zEILwRx+QjYaO/
QzYgT9IwGe+yoq+OoZ1LK+h+o8SvWlFo1lFZ2LYxKXmTSnttcvlWVGuXHCfLcmdevDVF3Knnb2q0
Qebmz4DAw1+60VfLRZNQZvfhFyitRToQWpwYFPihqphHe/zUYoZL5AVZi0C4LCio18v3nPp3u+K5
7Pliaj0lFyCrzwDVYvSAdxdUna/VPGiWuiPGcEe/wLTr6PZIYlKKfvMnV1IwGCUF+wUeOva335M9
1KaJ4mesquk9FDHjIbNUoCw4a0p650FA0dNipBz02pqqivGW3km6Vc/p+8ox/tJtq9R4WJPqURs8
wv9zTya18rvdKwqwH/ufQJFu3P77uu8ZVbiEhufl/iivfx7NcMvQUMOl/pwyRIrDLgamW3pSUaB/
ttMI0bDOYNDuciYfngpa5OcCZC9s+yRbBB+XX1mubLU+GBoa/xTAP0RLqH/n8P2Q1yATG7mHWMpv
jPnfZWIvTPLivouvAY7EPgEJ/PzaQi7pTmJAYKXvx0KTAOgIPFJrXPiitukwhZg4OVyhkjkX1jVZ
Cg+HVRzf3G+3fXdU8YRNL/+5fu0wgvSXBaY4cun2pSjZ0eHq/3iscE+H0bBgV5uCsyApRghAF5xa
ASRfj/Gd1ItM48PKR0ETDrQHZ2xsK40j7iiTQFkLsu8lua91bViwBAu6stYeMKJDRjkYhjSAk+UR
Nase4qE5CFax+wGdvneQaXBmW4DQGxL4a07CuYxAuXX/YnErgzTU/FK2gdEzxFPwstrhUYZGAPJe
jRzFXsXeA64q7VJO9h9n+4mpW5KMIdm8WX+TGSpVS1FRyVy1K0rtICCFLtZxstmbEm/PL4exN160
cXohEB/A7/p7HYkqjA4M+mDNuHCMhx0QyRnh01TnUG2YldaySQ1ERLkFxe3Lwjptlr95f5TIWrXt
ErsSPK7lX0A0tak2DMA9GXyYRuxEp2GnOU++NFwfE79bReTbhOYxzjR7Jleex9+C6+EYE5VZx0qm
U2bcSz0LJkW23fM8QlIO77G0QI23n8YfhtmTHfYIRkf3+F4NpFRBDapHroZRFQNsm4BOJrHvck+4
gSxoLiNVtTkiDkFFBf1Q3StSyVqzvhnAoLwLn1dj8h0fjtrjs8NdnVJxvh4Z8nIDzzQSUcPo/vHj
g/B84WzgMRE5FpPiJCWbKAzX4snTKt/s0t5z+2k5IPTUu3uRajghDqLGaQ0z2+mtP3KhDHR0rfY+
dOfs5x3KzzBCl9FmZX0yhsvuTMAKaXqIwLmuwKwt76ozDXYiZq9Sz/3WhHBYqsWo3pilUSxjTsVI
2QLZUk7dy/h+RgYL8OH8TED7W1Mrbk9tDWVoTDCi5ZTXW0NaBVT6LIamZsZqYGIg5lREEkgiaIHR
Gbhz8QDpL89uLEokSCLlpPSv5iU4x6wIYoaTQLjUHhpMouUBgr3lAftrxVAohLBmZyt/L0CbzRab
TyYN9Vskv+PBLBWKdmnvRSfbmKPG9WbEM6vh5bafhNy1x3V0pGieiGiBNav1M84Xp81TGBpZORBk
PTTvRi9PFOdPAHz6VpKHD7lJLdyuDnMIvaWiIHVub+8wk1lxuQfaVGUBNpVJANjL/0CW4a9tQF3y
Bsqvu6l3+qVVTcTgP3AYOkBNHMSmRHpU2oZsJFvplN13lYYP2vVeErKiTd4Q7SpQvX2To/uHIBnT
Uc4axIVVF+YLSh8jg9cfM7OWD+uZIhe8Y/UXpAen3BiWis65UWP8NmSC2EXhedvJnpPU6iWD7gDC
HYlLrMx7EV0Zy8mWYVlKDSimoZQOwK+RldT3FeVgW3tXHnVuLlkP2SiXm2oik7i/BrGy1FFNSJLc
Yd1WamJLFHXJIlQhDPcTLw6TcjbFqL7YRrjLb2bW5nrPMsAr62Lxzjq7idLG9OlJTEobK2bddBDf
FE9CFkrmw+nts702avSXtfsg2tlykEuc7wNS8Ip2yoKa4jDr8ULsAi2HxFqiYOwPXdyhwNXddyta
+UbTpiwDOMBW+Rign7m0FOW0RvjzfZRILhP2dLP/vQMy9W2fUVPr/pCLnofKRlHLpCB0ezT4jEnF
+srRbdCqRikuVZS0IOItxIFzoeFE+yIMZP5PIGTzmtMBYjzifwEyahpaJKyhyrFEdPqR/KTBvPux
NpZYKj4OziLHfbfuqHDhKtrq3Tm0jsvmIBof8w4ZwUZh5YTVr2FkJxWPyC+6VHtgUlm9i5+bFpmm
BewoIZr23WhKZS0Pe0aTPm/X5sGy2TEYcYtFgJ6BbXe3+i55wWQS7FY6ZoMhmeYfxTTZoFrxFR4s
vPO5e2tZjxDSscGDERxzioAuoCCICHHON5IkwQLDuGCow3RlOe+HqThEarOo4sQzWKhW+8rME3yB
H/HL51bM9zH1A3pm7GhH6WRwSOXk7nPcvMtrbeyM5+RVxVyaCy++MCkqF0yjRDo0etFQU50yxfY1
GtETpNLWD8iAugGO0MeksphBGhxjWbgbAxcLaHwFjiEKUzZtNcGR8BF2KEnXswSp8u0KycqBLQxP
hRF4oubnF7iLHb215kzm/d52du1uvgK81nuiaoyzrVzJDrZ/i7oPdv26IAutwL/20QNOr0/K5MPY
c0g4n54EPJtuP+NnQl3A/seXsZGUlsx6v8RIuHJsMx6kujbX1iYZZkJc0BycHUXbHuUuvuH5I1ty
kicer83ddA2/rPkhwsuTQEMfMbUge+pjZCYBkKQwZBJagtSwsq4PDjiIwntNaebOeeLXTlpQAeyD
q2vDSVmdtAJPaUkAoq+XjdhoexPyQOX+mKwKnGoV2mewDqdzRAtXCKqL5emViKH3N9zT2d6pMvsj
e/t8bClfA6azV++ovSdWNCWjeKF75BCVVJVHi0iKd7buPSJZcPdwgZ5wjjHCPOiWPO3MUPDz+k26
irw6u3BeyCa8kq9BYX7CmwbloWPN18N0TvZ5SghFD3A4ZFZf9kxg/0uDUPh+75UiGCfC5HpTxbHt
Jq1aEG4Mw2Wpa0sTnJ28+eaOaDUsu8XLhSzh79o8Rz6P0GwddNnoNhCNwddQ2igma4v0Ij/43NUH
z0/crAu67tZRBNWZ3pdCYYGFyLmL4S83nqgE5phe0nwQe8fEbTGBWkWZ2onCxmZ8ez00t2u3e6YI
q07W2Lj84F62/cGtDXL3EpiFSP1q90vAnUec94M1UsgEA+4BHPHVmwd+opyyGLIR+V1+VJOG+0ID
IyOAlvMWF8HM0M2j3tmWVm9BlA6YvUk6VdRWJNspKXKzrYLwOlXQNk2hq9oUBl/yiasqPPjtEQXc
ShRlTx7Wagva9m6NNNTrn7JPxPwOsqOqmZ01E7jbOBsHlhvqBIyMxOqefCrjspsTw4sgoN1QqIz2
m+GTh0h6ysj1VxmfWgZsBmd+kPpdC1vOl+ZQHcbxPXFyW9H5o90p9UnbpftUtH8MCf7YPZPqDJZ+
MHpVb9mXYNLVNx2i/ipQNqWatkR5qlgfOvCKEhNGNUKEngJxPNrqdDCwWz85QYBCn86E5TXbQES+
jnHCPei8LEDDgpuu0/rDLat1e+tlsYQSGdS/DgN6STeXqtbo2GuDtHhm8T6aLYql1vFZk32eI+4E
1ivObk5e93W9AobVvczCt/djf3TZMwPoAiMGyCHDT7PpKiL0yyySPqbMA9wRko0M/hqCBIuflsz7
j0qzYsDHLDov+1FctebHm1pWNpuvwCpEt1L+1nsbK5nZPnfwIKYdVULdPaw0RxhogDm1mICdOqk9
z1R8/ZgE0+jrtHzP/P/Ah/WKNc7YQben2kfCYfaiKEgY0be7T93L0fE3JMRgLfPIXjEco3sUn2BD
ZXArMlYrk1GhFo464dT9RLKxikrtkRsAyo3NBMDKSEWV+avonVS1OkYH25YqPlYbSSQLO1uAMeJ0
coeHvM9kjZJ5I5UmeVvfUmNFCRluccA2uRQWZRz1Jb69uzGaf5i8W/dWCow8qVGJ96sTeNig2Vop
g0qrAkWo+Y8WNYrBgnzxcmY7/O82Auy98O2WMVRqJ+gnamuUEdbhE0TfVQN9E3AP6Ly1B606AvY5
CS65obtLZpkPt5aMAUaa1ffp4mwh4GabOCnf2NM0a0ywoq+vadGERtWM0W8BB45UhYVBcEiBP4pI
j6n6NJ02nWcZy1o9aK8OCi0Dniq4gFeI8N9IFedf6X+zIrhPiGlGrK8V/S0wzbqffaZTS0FZbI6T
74lawoiUACbmsIM9xkR7MoWQiAQ8K+46qhO9uOcWlKodgF0dEmaWKfoyDEpVMUffYP4TMM0C3t7T
TOug0f0cRs1EWOi5qyTz8mwxl37VYBsi0cMPfVIPUpNN15hdkYDOGqrvbKszzOcqwdh21HhVz+8T
uw+PmUzQQ7SIo8xqHQLgF/0yqSJhUwa8TGYvXnd5RhcQ/XGZIubKjVqRVFYiWPasKCXXuf1cVtJS
4onbr/Hntm5huFvc1J5uMQ+eVwkucEB9/Z1A63YpjnBctlDXjM/T3qerktt6fCv57PM7S/PPBwut
CKu12eakNOf2V8BzGWAElSXjklEnWP9XMy+ALOv7xylt0eCF19uMxqJ6P6/yemNexzD7Tze7bqjc
sTar1V8tHhMKr6yVIMk9Q5rDrEEttDSYrfjW55073R7pl0NWTuXjGi482FSsQ00o3rnThN89X+iq
SSNOQQW/fFBBQvlozA/onq1pZWgXeJuK3+YwP1ATUxKJkdfazUBDyxvZJskC0Aeqltj1BpHT5pho
f51m97mT521dmWxUnOnJhJtBOrAWVri8yTnUhXREWOmDMkfctaViAk/ed7KgIDESCZNqWns976J5
GQwH5eEYSgjONyBHjE4Y8BetoD76L8EcpThvOhl7pgpi8jOJ8NBjDqsUDIcaq2HZ3LP158PC4Ew+
7wc/ENDwkHN5lszPq7UDnfuP6SIubUZ/BdZOY4mXtdG89dek1FwFrFrltNjp4IeSXdZJ45e4IkuI
6T2oEaG7kf0GKUTQ6vLidqiSsLw6xxGlTDpe86dFFgDzWfVPx2aRC22gZgZrjGm9o5PSdJ5Sgz23
Fq4UzPY1IwbignCcT9Gv15As6enp7Z5jHf3mgAHWsKbY+kwZdvyHY8OKx0OeREGRJqtAa26WP6NM
VpQYnpZJPji8uOBmaSw3b0ve/yMljz8FxurCEdsIICpr3kq07NiFfqWsalikqTsLRMEy+izsBzg8
AFFTJ73YWBsmX8HFhHNEqiUTUm34kFWI24/Mp4bOs/JJVMi1FrBDw9FackuEjAtMIQ6ERn3kcO/m
2ghKk99t93mnKd91JCZIhmnN5rU3n5ImdVHHrYzxZBVG/Bx2kvUFdNjrCBf49lHoICXuQ231bSSp
U2sXktUlfUu92s4B7XXrOBg/QxLPinFtPZrejxTS/4zft8TcZKi8deyKxi09rTWgHm67hr1KLs6M
obKouZPES+gLs6spKRxw6r62RL4ImIfiqeum/pL8OBlu1wkil5gKjSS6hM2nXoBeuGCA5EfymTFG
JeLbaEKivXIFSBQHlUEt+ZXIYDVcZsWHPu8Gsd2UKdutMAUM+E+NPPuMAgAC16hu2ekKowdEJJjg
ue3RdZx9J4ktwNNVHAmCz2zkzZTTdlaIjSgdKrv0BnIxA7aD2rC5Y6hFkf//YBszIh1bxseF0PQy
+KVcn6eJhe+kfkPYZmwEUxIY6UqjBlD3dro07+89xwar/eoGVqGTtjQp6Sa38R9Y73YQ92SjdNL7
H7mQQA8/2SxXub53AMR4RIX+loCd+B3EkcxY/7R7GLHJeQd8vSLg7Ejw/vrPYcn5ekPPT9H6/DyM
2rAF4iQgKakj5ClCX7c7QSommC57tStGfPqxSAJhf9GcY0I9lV87utsgxCK/zFCBO2yWxRTU4XSn
0s715vgfcb4ZYeG2yzssQnsPg6RN8/7tSbR1GAT7N+y68JQ41fjxVzPOwtNYnLuzQKqonXIKyV4f
deDyANTFCgyLSDufiFA0hognl53uimeVW2vDR/OInPbvmGVE0HF1EYuv8LXO8jiKA8UQ4em9KXBI
Czh4+arCNgPNmAm2QXZdLKH7BlrkiUzSrMrF8psrYufQ61R8HUrjmznk36JOrBMWgDEtout6bI+F
vFKDBy6mkA7ilgAAmOh445ibwl2zEj2bZqqsrjraJq5txfI9dqayGlVa9yL55FBSMcayccmrgzqK
W7pSz4WGv/BQAYzATUSyKjEO4hrX6iYPYjYQEDo25q9AgD0JACatmHR8l6QKOqs0pnK2GLp1ED3h
eHMlUDj3wUlqR2BEVL5IeYnnRJ9GAEiMT7GqZ6E3SHMdhEFLlmifCk/lDz/HfXf5U8tiGWIiyJm/
RHDIH0u234MzANaLOJtKaaKoU+udFPDcqit58TDPGmMdBDPitCysyzwjChd5FbgHLLbB8snIa0ib
IzHw9B2ciMdgRwwrUSIQ/zK9KwzL9ATsT2eYjpduy3lWHqHqk/gaPRrfTdaAvadXOTSE8TovAV6H
ealbLrQ2IqsO1V7059UgMzra6wtg9dMdwb/C8RMkcZWqyQXWhjobOZRbzYYbBrdrWbsk/X8htSzD
AwpuvE17VxAa67zeW9wHAU6pzULt1M+41fvi9rN2PbZG2s/307cHTyv3sdlCCVTaHSjgx0JXrxSe
fNHrQD/7OkH3d+ClINUGrlyTyaz8vy4qfqkq7x9Zv8JcMG5YSuCdja46IbDWRpok+j6gm7gzPROq
QvMpAfiUhfmBoAGZWrRWT6gBv57j8wCGYuYnXO/r/8Ut5ksnLdobWvK/CyfNq6aS+TV1szVqo7fI
V19T4eFaHvM3SUN77Ol+hMnkSDlCRlmuoABhLyh+hpyq9ZsIXe/kIX42FxrOgNH2a6f9GdcPRBcK
osh4lCE8IQM2IftN/sD0QWMh9ZtNnv3TgKAM8yYtM0D1NC4PtHDWUUrtIIPbR4kWz0rHKaTlxJmr
9C0ye82MK8BwyQa5HXXY6dI76E3X7s3ZdmrM46dkW0laSFPjP5zGsFYk95SxVX+axjTeJzEoSetR
GRRv79c3mP/HiMrU7ahNlJAO/dI0ypdLH8xwg0frIXWA3FOeNJFrsUoA34GLBxbEMrUB8A6Jlky3
Bs5N6uEQMs1a7g5rZJ/DlDGc89D5UM9lTIQe1dSkIj5iiH0WukZhMq6XhoOiGLoX4Ee/PrYTTOuP
utNG/lYUc0nis3tuEjwu3gz4RMQ4bSj6PqJcSMuGIX8hDVjZ3zSzbye2Olp4jXW4Dmylb9+UoEd9
J6zaEXQ9UYXZOLh3Zpm2z0cHAVUrzPYLfMTEcJA9YN4+kxMPhebLXupJNCbsq5Fsn4tj7N3ybJDn
P3bsQB8/uFSXcxDIlC/Y7rcymj+jgmeC4NU7Z18b+xoBQJpv4aLN6NPAyrz/Cj/WDGVa0kLWoxB1
nJk3EBFbqkvmkEm8mAXaMp6Ga+jQsb7LKyzcLhxSK1+TEVxtFNHL1i8rmPIO/MRmKEHAthUk8TVk
7dH2okhjY0hKQXUIfRR8xR/As7iw6VE4nvIKS1YfvcJsKEZz9lbnMFoT7UjbcDilDkdcDnuNDJQi
sH+OcQzgbp2OjKo56zVzAedXrqjvkdjnWhBwQnVOdXCrIUxlN8B/pdXYCarNolVpOcGbDBNM8h4O
JW0Pr9Fr7PkHpfK5W9+kcZYeVMfz1uiC7jCKBT2vZsrcFAmUgfh5Kh1l0jh/ie+jyla6mYCsn1wH
zS5IFHmcCX8GQDE+oSCJEtAzIuKVi6JUD4NvC5vSso1rSPGEDC1MGbPFeDZhQGRnxrcHKEQvbVus
wsBrBihQkDdHGJ9cwGP2E+v1S+TbTDr0KAhVT5lmoBi5I9MqsPO5lplerlA9AOlnToLRQ8kdjp/V
UhFFn3e86l9BHHnLDRBhGR7sjcxLet8DIAe88UVHK/yk90lLRt72mz9RkyB4lOBrQprz7c0KifMw
gW+XVrTE11ZEQiqUFxoKUqs1mR22oDq22cPBYI0SWXwdCrWCFP7lIt0ICBsT4aUZuNB67rOuovhE
zuYN8m5acXX1QzdgxoyV8yipVEGELhI2V4EknNX3f83bRuS1brMrIdMglhyU0ug4xP+/2ah+KEGq
kyqv3G3wy7ILI+kc/r94VWQ4XgXIoLpAiCUoHbx8tEoSiNz+REWzprmvCYHirElmS+NrgfLO3eNQ
XnTpPFrpyxlfwLIXtlq3z11MfVh27WuBJbxiMDN5aG5cL/SWywxtkVUm4pJgPH3otLhLAFlNPgJM
8DT5S06TyIeHHJpnB+gnWgaSVwDjDOkT8lhgxhToHAQsJpqgeuGs/9jz8ZmbX1nWLFzuZK1Gn1RS
SL8iy4GjnBhOThbjrOnDeKxl/s2S1eehGY0TDSdcOZ8HoKXVDunNbCjDbCNb4BXbCubbXvQLX1Hi
rbHNo+yhzdDZEK1BQC8ftyKt5LaVXOXUEg7/a+86b2dHDtGf0pqmO/7xL10+icHdokdJYdSjbxZX
ba9luO2XiEppJucSmt/fofz5ama5Odl8gioK9tc3gUGM3hsePyZGWfPhG9bNWTrtO3/h9F+Kwakg
HKkPIUosEdOX4pUrgB8aJYBmAw5NWABw2i7F8QZOqo1csiI0s0elABoHTblhaG9WK6ylcCyhRpgh
dhbmvFe+Ke+S4hj+lZPahXJqMpW9oE6Mj03wt81QoEFspr5w8P4Q7afOxR2JQh1OlNz8XLfAZbwh
KjweSOCGp5mDNsWX7sPAEx7fjNNo2B4mMuSB34TE/PUPSN3Yw3pk5EO9yVP4362KmCfyLAjwKH5x
/Vc5Ek28OzIK+W0SyZTIL+W10HMxxQ3vQRMlFTV76QYVdF9WMrOhLB+aOzSp29ioXUGsOYuCQ+aZ
k+WEVo8wsGonGpah+Cpn9fUb1pCJe07B34wtYzzm/JWUFQguMwC4vM+zQTiBE8WOEh/jcH1xfFsw
bcyb85OFJ32l/U1Y1YoOc0DGmErB0KnZjztMJhnFRt34tHlXMaSP8M2s5dHcLv6oupyVCYc7W8lV
7wHCOS3k9QBjghJv1Tr3IXXaqQuYtH3SNtHYh4smN9SayilaweE7nzKwOx+geYPm/MG7mF9cPogu
SR122eTan7tG1xvTrhB2n56YmruWTx/ZdoxqAAZfaxDAIaQx00kcm8GWXLIQWqZ54/5mVyNSzk6B
L4Z70cTyRSAYMwTNfM/az1en/n9TlwhUXd28V34myvFahhH9Om52X6433hUB+7Ly9czvNi9F4ymZ
9H24EEHFVchIKI7qRv6Hv4KEuJ64KwiR0OGejlpikwMDdQVFc3s62fpVECp4mv2uUAW3YgP7iTcJ
2m1Mn4/6LWuCQNvInFAEE5sGQEtWL6gWToExLrIJJLkoFGuJMhatUc3bmo4psGOIwrreKMB7VUdI
WuyQIvsQkl1LsDfve5KwaltPEAjJJXtvEQGVDfijChzX4QXZ/28vJVhpbfZ8NqVq0yvXLendr39h
U9I8YG00+if4bXUJut8VWXGle5KNMe7g1L6CDKULduxbYNxRMYpFhA+a1xKT3cvqUWVdseACie/x
4wN8roqHvbVj6GLBco6Pj2zr1aDHMn9DaXO5FzN0RHwD1o/dBNnYYW0H9/eiAa4f0Mm7fIYfVRaW
+ZHE8IujtG6T0HcewF800kT6wch0jgzVom+DhYr2Y3scwFyCkzpq5lc1HfPpT19Mw1qy09ahxsWU
vrKGTXIRTfrEjpl0vm9ZyK2FkawnlfKfpea4NuXmu223ocI83FL4fc24rECKqDhpAXoa+g29i9CM
zohTs/ZkA+Os9S/xJNf/YCe3eJ6R0oOf/6bfVf1hXBTx3ADgSVOAOVRWICKkO/L5nFaJzZNFQAzB
CLDXhegmloNMi13yzN/ymIhSfve02E1tT2cyYtmD6GLMu8PXVYx7Tk7HWnXmrQzX5N/5dXAJg4Ji
XIMrhD2+9ZAzsxOhB+D9ypbIFd18dWQOx0HpDVkDZXJhraYw6UkiHCmYU8JERfZsvzkSDBj/wwdT
G8y2FjsnFJruidVRiuYBcjtyUxQDUS24xlVxGvXBQ79Lw4fJqFl1PIXKS4asHOWHbeoJZUMqmnZO
szGmaJ+xKVvh4edu5EHo9yMZM+tNsiNXaGiVPxrM84K8942namHAqrqFlqtsOmRhVnDvbbJBq2V7
C94Hjv0NuepTGmHEikI3YNyMQk6JDAFE4U3csoTEDZgvGMFbxbUK/Ao8rZffchzuDM7wJFMxlt/F
IbS6k0ZOs0bNDYWK0pv++BjJEVqEnJ+ooTs7YvM4inNpZ7vj+viRVYHX87Opu+5+ZxxW+BmtnpEU
R0xzZMsJwiR4wjf9pyQEjpn8ulL6HqGHszBwPiNdvd2bLPTjdBo0cKfttFfoMYNDmB8ku2yhWoFp
ouHj8kWS6Yy7z8uncltl+m1QZTNmJ0wyrgtozqvJ6eRXLvFthdMBWGVeMxR0WBFhJ/irbW/cK+dN
uIvcKV+Fhm7smTEs3ZGNG/LEsiC0JplWgVRmFENopURfGuxlV4qwutnVo4Bfv+GgiCmxzMaM4r9H
OhNV82g8IRk0TV7tCP9PwxeOIztI/yWEFK3HRd0yjduG2OH19TTmeSmP46/pWa+aRu/QX51RykQV
Pd9yAO00Qlm2DG8uWZ0hpA0x5Ty/XGTlVuqMPikGDX1ye2mo0ZxXPHAcehYxt66zLsYGjkwQ6R4T
mmK8Xu5jzjGKo6j1Ac9xH32kprSe8RE/0BFU4X+ZxxS6YHeqZKHqKmYHPAmu5xmvRnm6w+emXmwg
tQfFrT7/NbX2RwN6iPzNKMjxkTMafmTxjwKRvOnXLq6HyXyf4pg/CfIMvEErCkAV5wLQNF3NSf8E
FhJcmsR+bkyboBU7yNiMeEs6XL9kaKgxmgglLdeqHymcl7ubCAhlNF9sbg0ssNLf0K0pfXSMfr22
mOMdeBLYHka4o545si64M9rYB0MTguKui7HryvBQPBxKPyKOEgp9o63nmueydXT/V3QjevHgm+0h
XblvSjI8teOvKHlBJ73J25TPrZs57Rta6TUZNO/xbPJzqCPdHj7ndviPylMPleDHHZ9cyiXBTCWq
5umbvrPG6jmBi5lfGeOiURUfC5RhG2qymSvWe59mWC42EKNJVL0hiCgSdl8CYCzegb3DWzfRW7vd
qAkscnHPI6eIKZ8M33r6w7rrI3dhPR9kUkwUakjl9gZNYrokgT5BbrDkrUfdxoDBVYx74fsBiuJ8
ErkQxweR9HPWTVNPQmgB6SA1zTb75v4wtosAIOf4/gh2/KTDzV0RIkszyMa1818fr8b+ZU8/Sj64
gHN7+sSWpWPPTwMpTEE+Mz0jLTAky1y47F25FosCartB64cP+suNWo1Enn3Q6OeX8kxQqv5xly6b
eqO5FiItq89iPoyFyYRLCFkKW/1T16wfvER9n9jDRv0htn4MTHHp6AKfamCPjIgjIwySkxZj6gbI
W2UrMIF++iQdK9/gR3K/PyovDga5vZO932X/b+2F4ydhR9euEVJIWcCQXynTsuofP9q6QsrvUF42
X5/allM7Q3yHk4Rpmhlw8+X+VyKIaMyaPipuFj/GULqssOOFLA/2kpbRZ6/wLCwWCH6sqTQHRx4K
yw1m/c0ObZ1SGvUYRp9WSTZPIdzfSUR/z2SQVGsZfl55KOe6Jf6AkmCJg+qT9fxuxZ590Mk9EYz2
waz99q/xH6ryv1qvTAt0sgzkRBOmOwFPoSywbWceejOTEzB9Rm4/xH6jaoQPPR7SUYtPl9r1t/A8
O4fxqmG7CJ9je01DkDiz7xbeynI6iHe3YXrbIVUFRYcAa3y30a218rIbISU0vOMZo5Avhu8z89Zg
JLIxVL6qwRmesC7doloKxuPaofJtKVxQQyDUcxZMqdSP4RE5rqVg2iwsyu9+FvBhjzAPLzELO45l
39XpnXIMskO1zD15s21TQ/hb/52DhEsUt8qsVokhmRuzGJerDI9gySmnyZrhfo+MHBaBJv0GnsGR
TFBAo34PoTfJmdIFDFFuKqctskPQ08QgKA2OVpT29YNfYDKbmAgqcnyXRxFQtEq771VvP/+KHbCW
iwsn0trHBjVuwEucE9ZtlKHPZZBczJZ5/Ssi/TEv+KafW9Y81/V5srdFB2H/omtNgQKKUDsHF3iH
kYIWpSie6sIm1QlW3xkzY+M1wHWYXXv0opxxhrm92UlKX/kijvquKVm3uFb7SXu038V6oHLMXAvs
NwRtB5OdGRXKfKzsC/zcczNy+bplk6FMK2oQReoH/To3HumHth8o2+GwhkZQyl7MQsUzDU78HSsH
Ikmo3pKAqwAdTg2vd4Dhpovp5lP8uwMDXr33OLMnc695TqUvZ2NDA0QKV734hNs6VZKSOdjJLc8h
dAyqRw03in0mhrNWnKuSrcpvopknKG94V7cn31iqrXqNneTnvvN+r/kQwJTnJyGMLqdeGyjcFs+N
MHvJDt0dLu17oLNkBuwvUViYeIpv4FVjVTdRFLAC9URmzakHo+Sj0DfaSnPphls1NTiV6vRRLIlk
e4+DjoP40F9JVzSSusFO4FoQIxThXq2zvuv/CR++Q/UaeO+/7BQUSDxSJnnOQw0nvdjYSe+CUDjd
NsmeDiheZqPzdg7jwEumMHG83cWRe/AzM8T0nXrMbNTOKVMUH4sbIa5rRmJufrygZhBy9xQUQY8t
61yZY14g5ltDgGNNMJkObCOoFUYFdQR5KvZpP/GbXiuHNLWBzNYOmlQYxfVFBgCNDz5r5W30tCgq
AgokqKWgbeb2L5S3F2TUS5D3XykBPTRwdLQ3FTDZngpgatFtZga5xWHQe/q4uhefC34CxZsacsvi
djtxCNU4nnRB5E3ib4HXRvwFZV3p1dO060RNbP6edhhk75cojyDJeo6DK+M2MTQwtWBRxMKDWDBh
8cNtiIXa8ZHPst+5W2tzRLmifXIYixXq717sgfUOkxVLA02QY7ucaGj4lTW0ao/6Aoz1BPryjj7M
FyrwfdbRwIagWmBQbHYgOuwOeTaI9zLLBSGGii4ua+1IfXSB/X9HbC4zUkBWkDsY7uZrBzClNq8M
psT+phPgnWQZuWZyfDscSBUqrVQHNJJxse9u7wJpRbJ6Nm9Q0ra2VwS7lMol0RTUEEJqWJaLI0eJ
ZqstjCUr6MhnS8wYk/siAkMgiUdtqLZjFuvJKEJDEgmyXcAYAoMYDhAsKynw1XWzcXvuDR3o/5QN
u43CF3Wzbdwql94onqPStU16r77ZMUl+5ntehoGSuE0MuEfAPsO9+WdomgU1I6EyNDymjuWvqqAC
+9CFzz/2XyAn8MdnSSXD/HrrYiqbH3j42sjOO4WgBPwmw8lqjmat3VML4HAHxmOUQMARzq8oXjDd
DPUPhzjdvMxNbk5AFqR5Htj2Q8EIm9EHR+Qnbq+ECZRjOIzLNgLKBy71WksM4v5X0tAUyNCg0g5C
itIuwMvHYqTukMfd1XB4ctqVDRh1+0qLR0Z3pjNeIKiNcDxkMskBTIBCfCdWA6wfQ+mq4ohHhnEX
vK0zdpUWE9menyfyhi/dM/QS31+dbVAbAKvYtGts4Juxoq+4CHM3DygqX1LsXuZIvVLJbmO1Um7U
Gu6u2gckJBIfZ13vMffrhuuyOik2Gpa8VbS6eDyjNKEwLsJ0ApjN/+8KIEz2SkNDsaejS+uf1RQE
s9IXy/fkQfSpZAS3F5Chzh3eqvfUBLJ03iHUkmr+Xxk5AbYYhKjYiQFOInGthYUvSmTJf3cmwChc
U0Az/0SWjb++Ui9zS7MMNiU7z4yaokydwYWAHa56eToisBQJBrjvjQ3u4QPYO4eP0nA1DQpk/ajp
rCyxG+NaO3LVqy6fazUJTpdnFFjCZEG/ISz7a/EkbwuLA11m0uA0oo494kwsGBqYUQvWjnc+x2gr
VIdSmAZlAdCeXSNJqkfRjCK4PJ0l0YL0bcOvnG0nj8MEZvXxK0cjJ4ZkREjOT6IBuT2ySTCP7hI8
SpMzLUvKzMfaiyn+1lbVe5sSsex9XlU4OYrgnxl5co3ojMCRcMn7xYkUcfEg3OJiFPpE/J5ZcOIK
wXpAhUuCW/nEn6RnYnRMGXCM7k+QYXQbwGkNgmpg40NPOmw/YwRoQivRg1CAH5FW6lld8vlntBip
3ta2IbTGBFIO1khkf2HE7n17fRVq/wjARVOBe9FukOjSjLrOCasLWUIlYNs3Tav46e5UaVGiaC30
vPVN+M8EiHBRylNXHH6e14zFyH60Knq3V9raW1EBMlaD0c6QwRCR1e7Q1lZDAnoqint4JZ4tIZKX
4m3xX4CWhZk/nSrKFdc6Llqad5WJ8Mx0wBXQPuL72jQ3y8eIiayPS4Q8xHids+aK2uSv/KaDXuBH
OhqKMoFVppVbd4+jllQwcCWuwenuZDYY1/j1kdlWl2r2kLF6yjSSnsRK85DjccVjKMVrikXUOvqb
BOMSjf+7C/lLhSU1JNr3IwVByLCPoCG3rKxhsW+MHn81309YRpLperbSD+2hZSQmR3yz860CwQk0
yUpiaLcc29jlPq+sz+wISghRzsP7PqOe1bN5OWQBESgzt1TTXgqNFzDyaXq+dNgi7KYGxoXg0n1v
8dae3FMuy/m7bnJGSrpVkgfphbksy0GQGJWOdxeYJX7RdUhxlshlp8oVt9BCAvFiFhiY5bDJ2oo9
NhX40F8qoRaCyMmBRUOK+JbZkn2jIC3sicSMIrplWh6tctYh37OKUwymc1oWt/lN5F8qkIksoPOS
BeYUu7DuxFO91kG9ciltsH8nVMlHB0U6IOc/XZeOTbEFkZjPs4g4vhcYp7g+bIIudNnmd1/RYoE+
amIyd7rtiOsyAVuyJ88/9yY3e3CNJD3cN7d/diPJsizPCe392E9y8FV2JjPMPn2sApjt7bpa2y1e
PebZr4saRq7lW20bMTalbS/bpQKsthz2kgHUIHnHb3v2JQI67yMiCHmXXRv+AdBLEitTZ2U7TbW0
DE2qf/1J/yoXUDdsTegSUGOtnHefw5xNa+DPv/EXQHLd8+lKgEaLqheJdGjxMzzusNQ/hl6kehnR
yx8Oc72i+/cen+vorCsllyPiCzWmR1Sd2KoLkXw5fQapBp4+c4HvmtxHhlDpP23e0TXFgH0P/SYg
PI+yjaqtudJLiqZS5QYfBdT0WhQUctA9JoApuqtBbfjnD3S2wh6g/tkSmX9fBaBP0wcQDxJL7WOS
Aip/iHlB0iYvRXlpTxsOuItRDu441W0i8bW2KjZO4ylUWlKe1FypkerAZ55nfinLUfcUJ/u+8h3b
NhWeCjSTrrS/ff9pp/kQ+Cp7V0nI8ILHZU3/ED8FBvhpolKtFJqUsPrGfmMcmtsI6FcA10Q4eu3X
F0wNtGA39goCTxQFYrzInYU9YQtv6ZrSrubigvz3R/rFJ0FNnJ1yZwBYCO5Hn4Xfa6woilWF82vR
7yRfWs80dNnCZd/mVuaZ3Pn2ZJ2FkQ0x9NNaFuNHyA8HmPJbD98vssebT+pS7/e2Rax7DqGl3u/u
y+PtEVuJxNFCmbN76J8pYh9xoKkX7eMU+K/+hrsNShi4DHeF+NNkpb89rt3Lhg+JP3+q8hhmT/if
Fouq7z6/MLk+qd7PnYr+8uvQdLe5WVwoXr2EP+OnsiO9fBGZBdgJuLmo4avV0hrmxj9x42P5RcpF
QI30XjNEKi/+AXaV+wULeQFfny2yl2qIih4PGg8gM/wbxP9EUk6fBoqxK3aT+wdZXeTl7EAuWuIL
RUFz0V592EiHA/6bcP7Yxdwi3JphUizE0UKG2d93cv5PVnUv6UNkIOAkR+HXh1ok5z7ASNu2iZFF
oyh72Xql6V33ZhFFvyfDDURrv884bOrapkJqT1OZsIwwP+N/946QvBrPap0iuRi/WoWGWFIatFuf
P/+0PaVPKcbYFI7OXADQYBgbj72pDv4JNB72CIqOtm0OoI5k/f8YOHZrUTwalTsxbLNP77ligRyL
Brm/7ssUGhZKWaMhGM5D0yy4cRf79oK9Qx9P6VImh5NpYUv8VtzsEHyutH0EMMi+puLlWGD8hMAw
dZDBhMl+yvig8tINzUm0BEXf8uTRbd4RAg1gEeVNIndWDwpRxWjuqvZRwWCx01J7rGWmeWrMvj8p
kdAsqscpH3Vmhd6mBMGI6IpCFOt2WtRPFUx//atxYrEogWxHifd/ejEDJ8y1VhoqLdLmWi3AFXY3
UIVjwrNA8OIAbHlILBzo+2E5rXg0aVBAtW0BBNlBr8Cnum11DhA8YGC8Zu8w1kHepxN3sfDQVRmV
q8OsHSzwPB+sIks7aqn7VDn1dhv5mpWlXNIHelq8wpsaDhxJB1LrhgHOAhRYnaHKalG3+C9Bu1RI
g19KslhLPIGB6/6q9GmeOXqeYJJXPbSh9ZxgS0Vmo2arC6zE48Wn1tOoDkyZF68F2+7l7ywwntfd
jGcpSdeTx7gzAB7rgNBMNKXOIWQ1de2m4FyqigC4tWXaO7CwCnlDIRWQpUQiMlSog8a6nxvDUnp2
/qJColaYDwrxlxY/+fEnK6SwDSdsracPnCfyhwHcOyzTIdJUF4RD/mczRSMJtVA5Yccr2cbuUd8G
8myUamDdwsMSHfbw6aGjBz9qB5g4Oj1rnxoi6QAavt0Ji4LxX0zy5CTgP3Gv9gzo+ESV1xbnxOSu
ZLkUXT5HhzLBhmOFyNTzERutuIrP8Lp4puQtDImCDM3AWE1ObGbCVMCiX+4VydVA56OIBs11J45u
9TDdhhsrI9gQ18/WyyFzBK4tTcRLZako/znhUR1axElklXFe/RMJxwq1FUtseUCL/hFXRjPmVtN2
wr2EsqzH/s3isjy66ZqPl4DC2mg0MC0ZHn5QDbQxNi5FFgrOFT70q2qKqfO6s8vABiCFZkL/oIhT
xnfNHlLjgpjcX/Skm1ZOlxR4IdLs9ewmN7KmVQqTdXksCNYD/tuqBR40xKKmB8O5xzik7miuqfWX
8xPpGvkduxMqioyI1aS3KpiFRl0a89QtmSwGJVNV9ccWf/xreCevcOh4udA3MeEEwQEw9wsuFxyi
Ni1Qn0N1PHdoDQTpe4vj6Hnxa+YKllrchxMK1qJvKqQiys7DSweqi/1pFPfrmA1atZ7h6J/8A58w
t/qMXkeXWjM07Z7SfcoxN2hlBCnLBfCTd+OuUIdZMFzwcf/WFCSamFm15NcTMSfesg+IUV4Xdk4R
XvUQQufSqa6zqNQBkVn90iZf15FHMZaMQ34cJjCpzEYtO9jppzebUC9qt+2qc/6T4n8tNZRxXZ0F
OIIXLP22fF5bY9U8J/hl1YURh1pwq62H8iDluh6Y5brXbUYhhh7sna6DOS5jRAM1+VSZOdRDxu8r
NSuGAIp82X+XD15A/z0tZdXAuBDZP+g6Tqny2eni7gh272B0ZOs1CEGH2HapKx/PdDqCKp0wGVrM
+ZmIaQS3w0CdUD8I7LnzWR0jHeh5M5j3rGW5GRskXnmJtDTiaIcb9B/otV4R26PRpyekZ6eBnZzB
npIL+jIvdlWUZyzTBTqn9SATLLjGeWkJmSbfPR4SLiLVtBBAszoJoFlV8OHCE1gq8SRvafXdKYKm
fIP0xKzBnIN1vuAN5hjGGsItT6beE1b1jb4Lj59N9xehdIAMdZx3a/H4fBaCYmw4b4OHlBTZMiWg
Imo5IG8Tu0oSgCBM8iMIzFEmlZc4ZMMn06J8f/eticRFtpI7ukM8flvqICIjhiumbGsed4Wrde9n
qP4P+H0uIbWIf0KKVN45lUSPROrDZI8AVn4RHMXNZ2OXFSQfEbBUzAs903z9TMdTlfHu0CyZGxeF
lkYuh1hddR63Ydn1eBD6ASqGHQeClbSCJHBosTI0PrrcZNAU+4DzZ0Bbx87tvVHw3aLF0dBDEERg
uSCtLXXS62gy/NTx3deXkL/6vQZsH9rJeC8oRhzbTGjlQVKg4IH8L2MwF8gxWI3Q4zpf7xOYNwxH
aIMr3Blu5R7GUYqnpHGdeCh/toCAJMaAcc6cDnhUN1tqvy9hzTNlBMgpPrrfvkKGgT8CsYkt466r
oramkQRSBC9miyVOGhvCkW5NlAoC41xYyraZ8cHsJ8S3Z3uU8TWBVBOIRuTTZ+f5py6GRIA0hS1Q
R7zTC06Dr9wxTUYS2bC4vXkqL4ckgcRi+wmeyHbADiEFD35oWgYukAwdmSm03Le5Bs9XMIEiT/l0
Oc6V6hV5+skGM2z/B+AEnGSM89T6PHCwLlip0z1uEsG7e6C11KTniBjnf845rBrfcCzoU9bVyCP7
UadHIhKN99stmuGe1tPczeM/SSP7O7vag8MRUjRx4iLSop84S5SjijYDMTvthqby9Oglpay7xHoP
FF1kiDqvfb2aOWQHeioBq+lfPHYnKfCxN1zt2QS0z1SSEj01mTZwNyvj57sTltOi2GCRPqWk1zNt
im3oKh+VY3KYpEcJl4KPLITGZ9bABvzpao/kvIRIa8ho0mumLH6oi0ggePaoVkQDGVTqAiyeNpmE
iLzNLG10gpCjODlxKG2W/g3+x36SXI2zYRDR6YOxP4nYRaKD1AGVWxW/5eX+jSMHaLDPdrzu6eX8
6D8Ir1tCHC6ZelftvxpPlqSGI+V+yjzXKuTpBFc7c1OcVD0j4p3LPEwDTgmaAwnVTGC/r7YXPyCa
i1fZ4e5CIIufqXR8yx84LQXcJalKGBYgDzdaxA+dX9f08oe9RY0xAt0+tnix9m6eqhTnXGd0cHA2
/Qr9OMfMauVcyx6HWhZl6LJdt7KZv4DFGk+UclsZX2XlC0czWgx9OTd6McfxjB+u9hbe/euhYP/X
wrOyTCTBUnNL17N1NC0DarkMTh/DjrSXJlIuwjeSKnLtsbO4VqIb6Wq/4Fi4/R9tQaAFVhhetisg
rGebk3CXpybv3Mkf/Bg6ZmfQtYGlGE8QNa+7DFMshR6UDhklkWJ5lH8IF17mDKcj6h0CLZ3AEsVN
jkXhMyx277pbuHq/cDNF+Isv00p41pXA8OZqpEvhZFw7flIkTcfWW77bkOG6bKIWO1j8F0Ukndc9
JdRdhUb7WWHHHY3+LBR0fNL2n/LsavUlkUVrQXbkMMPIv+bf5jXIW9nNGuuIg7QBe4gJVJ49Rai7
3jLIwmDygmvSjx1j61U4NpGeG1PzXxdzADC4999a9RDzpieVuA4wKlSjeBoQLnluWk7v25sbYkef
DSpwFXHo9d9iRIHcGcMksUOPH09akHfzD56Soc015gyTM2l09k0JC5K7XuhEbsXw/pmnAFNBQ+uh
JD4tp/SCfA/6V+lfzhFNUxDGp+zYxApysduRJPFNv8XnL5EEitqufJiXcBPEUqw1VCbl1fLFW/nE
z5tSsVux/OHKms8nlHidw/lcbpbteLUgwJcFzf7mED93LZmW2LOTGUgfq2E6EP/nufE4zzhLX275
IwJbSOAxvvJMgZFHe53g9pozATooY0R1WvGSWdaEtoL1ZsNg182DFQRK3tci+mF3Kl2eVJ+c33Yr
mQCsVgU47x+pivBv405Oc+x94jW16GrhpUOqkztMZV9/IQPgOpTUAInZn70TTiOFEMA8ydCK1Cja
9eo9YeHP/x44fYvUGKh5mTRqF8TJodztuhcv8/g5AfLABkV/4b+ZFBDEoW3n5nr6M1p3TgKsrZDs
DWxj1C884M9CLompcpugELTfCMadGgndSv7B1rf3Xqf5aPXdZrDxqZDcp9WMnQj8ojLquDaxO7GD
OJSoIZeSjSrTACiOnbFbRMDcuWzu7c1maybz+ByvG2w7IAsB/yi7p2U04apst0z5LR1uhMvPXO0p
fjenvGo4vQzZIOc6eoQGvcGRrGvJyCexUcPlGAX/rHLz6Q62IN9h/X7z0QvLLGHhFqixdWZOasAq
8huU4G+ojOtFyXydWTqBhFfin0Uy9wV/TeqtsDdabgMNw185W/M+3QmIrI6RgwbgtsUj/+Tbe21P
1xjJWtuBaRXmJna523JdvNff59FdFDKWAg6SyYtAjOo71i7ozq1VzSYOJJ7pVGDo6tkzJV0zU4WD
cYNV6vnlBBpAKYcP6Wl+QQB6JTyuPViIVip3/ESNUIvT4ZTkiBPiF6pj9QtVpA3r/pv1aVRrbWFi
1MWzgdIzqsp2LOupVcxsgrueiFc9nmWWs1itriVf7NRt17y0qvF+YQW5Xi95HtEGgeo3iRstXkCH
c6TLl6GhcBvH1n8e+PzmebXURzfeUtD5C5PGrskSTL99e43G4lTTwp3JbrINvi8Xo6tFl6QnH0fO
eCgLjgShP80HQAnxdKQ0TsQiaSRH3cNMZhpJ/gvt226CDZvnPpVIAO1wIxWSbkv+sXr6LoSB9POz
2cfQY6a1+uglNRuRbKielnGFJmBFifZFZvHqLoIgKRSSVT+F9k8GniUWBPol8GOXLV9cn0a4K3TJ
0XlYXwF8IDBwpRwzj5Fs+u177qmRFaiXNzqI810vpLlfieXKWx3+/U4J/bMPTK5GgrqKp4TuIdK1
hIEuUb0wveab7Y90COVtdbof39PHZ8Fmy7oq1CJJsJIr6mDmy7uBxrFQHOWxdnRoDtzXrM7iLHhO
B4hlAFkdZKK261Agio43wTNbMY3wUuT9oSBWrwed5BE6UP4mXkfcGaB6TIPWDuHbgHUvjlju16ub
smHkLWJTLpjnsU1m9s17rmcBn2Pblo0Ovfw2U6YOCMqH/Jp1SsJ3Q/VlJXUK4sVgtii6ibKHsirv
bWn5jN0wp09qG+P1HmpHpvYb+Bk8yCXVEcNlNy3QRONdfX+YVJ6SQBsjl0hllSqMRUrt0ylIHsm+
7QMCj+ZCYlBw5vE91CreF8P5UM3nftRWoYGodF2+YJ6sOSWBxgjjGIkyTyswQL5hjwmBsD4v2XhC
P6yTac74wm7fgSvrYnKENJZGJz7qFGp8cSxLBxGmgfhWH1xMueSPzr5wIqZH+/SrBLqbbK9/AClU
F0AxO7Pf38pOFw53U4zKVllgj8S/DrYA4y19Z29rJuUGXSpH2uo0NefAP1ZWFzf8BztCg7e+RbnA
Nr1bSI8HSuzRr9h92Tt1pF8AT8h62a9ycMhX4TDqilQrp5YNn2qbLD4bG2yJ6i402ixC3rTbRbEp
qdUsl4CmgUxa4WhauPq4xQlERbso/tNNaYpdUkFE+5Cr2cWgeXPjdkCaOXsarwuLchi5Di68sfsy
/ARwLFOZLYkf2S719Ev0xHr7WkRchOd1lv7QNVLu5/3Vs6BZyUC22C/j1Qw96SMi4g2n+edxHoXu
8p7aE2Rc73e9IoE0H4z4IIc/RQIvpwfwb5AmfLbw2ffl2Kl0XIXs6R4F2yM7LdvEIxLFsDfnIQ0J
sEd3trapbA6OYUOBWJVMPE6JFjO/W+rK6R/84UODUoS8b0hoTM3Wgd0WfyMfTC+l6Ogq98+AM013
F+jVFAZvIcHiNyq0t+nxEgc4EXTPPd+/2OVKB8oOqpf89o8JA+Yo/u7fchMfyNvtnUPWblll5Ozf
s0L8YtheWHDA0SRDXpgB5qfy1GTPu5u0fd/6Fi6emCLA7qCCR5hcjlQGRZz3m8OE3xY7sqZMoAdY
e0fKsMPJiw7al5YZTf85qzOZrvnAebI/RzBodrtSapT2dgqNMc+J7Md1oDNqRz1gtg/cymwBbkc7
orTR/jQ4mgcJo3D/Y/ZSvZmyZ+5gqTojqbLWeHTgL5mXdkDivGlJtBraC5CD8t9EDCLRYpNm1nw2
3nQZou/PEHF8EFsB52PrXeXnjvRK7qAY243ceajRdGvk+3e8s788XXPgzppck14lTjE3goLpzK7A
WjbqtPkb8SHoOXayK2mhLHK+fZC8/3H7dMZqSpC2gtroINLTs3WJbqcJxHUBPeoDZru66QCQBRH+
bV2jsYlpcBWQ9gVB2JbBkXGHFWWN6BAECTw6GjdHrGYF9STHy7/oufNf3JhzQnK4b/F/BphM67G7
Mn/O/bjToQeTypvux83VoKNYTZFgLdKkE2Jj1l5Yhl1h/nBqdBlzTsTuelNggJMwctXK/TBonTMF
4wKNWIbGcPAfBqCxrpfLwShXGLhJu119MDkzvFu0v+WgzGIHSwgZRUCP47xFsirzWXXOG2bMLL+r
YJEoAXAodY8vKmMZrmNCDEImDA40MTnmyRqMIdwVVL6ivOgUNYt72u/hGBB1rlafsz2+X7c53RLS
XgQynLhNXch4KPSQQe0PzXrDAIsumkAImPWEqQju6vGzJKKb456SIgCWegrW2hRHSBGmOZVlPWaT
nx50ixEiX1C8axM7ftr6JohzscfNBymuGlvZsSZNbhDE9giPXa9/Afjs/B2C2U1M5+FY42UpOea6
e13mPrK1Ufi3VSKiUbuZ8E2MR71WBao18W3YeKQffFkFCCod6C+TIDne3vz9VbeWjBMKseWtD/4L
1BhywWnyku9lQS8iN8s2H5wTvCIER9dd/g8qobOPAXGzi2L5n6Niw/tfDGnCNJmYo68Cx5A0FIYI
nahvbj7skA5B6zre5YpWqNeRvk9OVsbPMATmIfW6+pyr84dMJf+RtePoVB8FuQr2iUPSzEJ/I+Ks
plQMtGRQvGvMJvL3CYFfJUp6G6wkaPu1L4MI89T6WaEi1PEvYCnhoYtwN8ouUBPNF3JIuMUIAgMY
i2u62nzHL8PjwrHyHT5ECVFIzXrGkKbKumJ7LXjMMEAPAxBmCdRJnpUTObw2O/Yf22wbHH7DRPO+
dRSrugMDjQV6g0qq4pWQoZVRZJOBPlyuT22lCLK8yivqMWenSdmBpQQX8X4f9Tx9ydiuwX+CUPbe
XR26Nzx/cukMJpFAJIAYrP5e4vCgDTM+th7rn4KH+nUaWxwvGvQ9v0sRPwzhpuO9BQZM7Qcg8K+B
FwpNnv7R8kc16nc5p8JHUC0XGbSNaj2TWW6Vx74PFKdsu0MT356rLq+1/XshKrxEoITYN2A64GS5
qpB89jIChm0OW782GszyGAwXMm+6dLT9sFVQImYQ2AX4vn1khhKUso3j3ROqJeT5wosusLDhN1ZT
GUxYPQmf5DdttgLXq0hK5JRPS8g10aVm7bZTCm4WRcbC83PkBMeJbCnfWEzqfbN3LvNoLIc7yA15
C2ijebGEFw1Yxx6zcUNmiOrGsgN9pvDTIcV5ldPI+951bvqUVY0DuikwMomqk3jtP33Pmai50pOU
yNPefOETfzOEV0frnRL3F7x8L4eQcoPIfDJAnvHukEq+OFbqEYvPZCUjPAI7q+MPUED0DQm6bBV2
RBb75Y3a76UDQcnAtZE83x8k31Un7kcAhKGP3eRNdWiOlvI4gpJ10PRfGV4dXyDG39VIZebq/9as
1bVpI8k8yaARPjxRqm6ngqlYnTfeYI7A/SNjoUD91me9GR+Pg76HD33+V+sGHEHMHRsaAX6W8jvQ
lwevUAAbMZgzvVR9Ck5lk8np0uch56DYokBQqcIy8cBBkQf2W/1TAO8KqkYL93Lc79a7BXLZ6DR3
KHgVc8IKpiFJgarX9uUNp/wg7Rhe2zlDHunrCMIeZqkh+SnIWPMfZGoyTRaJqxAz3DRUz5lxa+8d
exJZ5Li4qL1Lhvu+8moYmjigb/2JehjUFyQ386i/2EVvHyVoDKyXQE1zH9+m+ybT4ZwHwBEAnkkk
eh7B6250aMlgAVFtuG7Kxw6nnj6l8oWsgu7KSdamRwtQA75Xwfe6TNfWp0rXnVw8kXVy0zAEANoA
I4dWLdmnVTDJbDcISejLnQp0Pt3Y5uni0skUpxy0QEvPwA4SjQGwBqrQHrSBHevEVbicQzk8hPxG
qoaC7X+is2euTrA6bfy9aEh8aUc8ZH1OCR8M6SLwY7wBym0wzpoxyfHfZHgSxMQhYA2H26McDJ/5
Dm9I8pEEG+O9Pi8K81pBHHcRaf8hmM9AfcaNiAZIVCaM/yHl4vlouAv944jxa5gcXJi4KGEGreEI
zadRqtWRHk4c4J5S8+WglL3PnVCa8ajn90cwdGUe33NYtLdoFcAKV3SDr/wbuZi7tqwcdg4hCZkg
z21OAAtAMSe+QVCyJ+HFVSAXIBxgJiCWCVoFGS4DtJHo3IHiVnXRhFA/KLotOwZyQ5sA6iWiBt66
FPWzwjJ6xc/5HX4diAgq5DkDhTZl2NchqUbHFwFbrYhUBTRTRwGQQ8d1uDMX1yG9H3zhU7wbALTf
JlY3vUVEfFh2s1SkSR/ebqq4sY8JCImSjZ8NIFGHwnx3E3zfih6fXbs4Qm/YuUq0CvYwGKDAwoXA
a946V/Ossj/MH2DJxbMGEPxferJtILhExlG83R2s7sRjqGRN9mfCpuxmC2kFFx7wWhItTJe4vf8P
0KxJSR0iGnZe9O6jEeA8x4PM48RoqPiA+cmOUT92hy6WXMHuSfeDxbzPK2yiDF+50s/vQPOCdZeb
Xt833CN01UuLVxtzxvAMPityoSzY9DqzKUgIPERHbv/r0Uyl+S8xZwqE+4LAzupxPThP5mMQaR6A
gBRH9GZuRbd7CL84mkHQwEn0g4ZsPtOnC2HVMuc5oXidrYOrqzW98IIP8qqozqtyx+48L1jQoBHe
j7QUVxiE1SckMqebZLHGpFCBC8A5V6ZAMnwnzn9sH1NZwbFBalGqOdYEpAqFql2Jn8G5/EQICWS+
ytQ2kZQttfvkcYddSJr+cz0zSO/gMvhVqLGblJXHzjDHhMV/+1L47Hvt39gbvJKOZp1CmGoM5J2O
TisvUdx6qfCpoXEr+bm8zN16MEDpXPBLmJZGwzWYPHYcRz5KxIpUVQdsC4IKuxYunoLhgqCVzCiZ
uTpPdJ16BhbUPneDzVxFUhWrOY3/qdaqj8NYycI4GWVdUet8KZauOlTqxb+48UHc2+ySQy1NVzRU
ZMDt+pmSqI0EA0nDteX+ofVFvZ1vl33hIIwa3weaOHisAhvcoACBQsqWqnsPScz9u3NBACuq2izF
LLzL/u+90UnC8puQ0JGpIUG+pfvnGy4Q6MPMt0t1BDx3UnEvvQsn6c1z6+8JIY4X9xtwLq8LE9kV
jA1oA6tdzJIYG6oLaMTrncKB3ElVV44QELstbv546s3ay7iHbYS5ocOKZV7Af1FAp9eY3nLIoBKm
J2DJgdbp0HrrfdEPgBPtVEMFmBaIwTVRxQC2FKzAeBcVyBMZdmxuLBxouuqjXraSBgAyhff8L7xZ
mxlS/55Gjkj8zyGzLcRrbJR/Xv2XaooSso61pTD5YfCyW9/VaHOtkIXqVWEanIC7yFK4E83BpGHW
TUBMAp4yK4zjcpHwwUfzkeryIPh8rhCwNkN5vx58qkfF4qhjgBDfpTpS5P28CKRGf+VeuguLKY6x
CBMOZsk/sh9JisJuuqyujJmE3fSw1S8LFRstPyAyacmhbZfOJZsuvTF1iIx+86lnSgNOJzYQcqjY
40L5fcfvKj7YdqdSa2ohgd2vXYGiLNm9q7TebeBeKAz+zIySlPNww66UjqoBXhTCKfi3ywe1VdNt
A42/k9IeHFAu0cQbirRxbkvufiNJ2Ka4Wilj8IAsV0kE5Yjrst35o2T1GThUP3RM1R9rIKsfJUMN
VUp4tLYT2AE+6IkyGqB3UpsIvXGzmm6lGaPYbdk5ngLuQdj2s66x8VbEjXbpo/3b+7VMfQbwrEXF
qcFFron1X5XzoOWbhaDv4U1uO/5xpJMu5+DO2te6kcjhsHhUhKCr17sO4NTZSyH4YtSKkJl5eckB
65zO3IrfbUW1pBj4Rqe7a5m9IapFOw7pRqjWJFm1wJxis+b0EgQXgHPNdcDRO8QIPrrid8gvOGQC
vx1EvaasSh40B7rXPfAb7qVkJuCzWDiu641VXyVnkp3y2dQ+YBbWb7/BTngJkklaaoKqHHNbcz8p
8HgAicdewGhc8UHxyt37KRgTdaBpYL3bA2B2tIF723B0j6YKDHlvkfKitkeZOvO613CK3IieKN0f
Dr7BAH819HeXwn6NS0ycmZhpQ/Pl7wpbwAJPMdu60thjmW0V9sbtLf6Ldo5cXotwrJV2COdaDm8M
O6Kx9VnLlOwLbpQ+kIud49I3dznppdD5IwDlppfdkjURHCN75ZCVKAQm0PJ5vsEdk2Tq/ck9wILQ
U5hDh/i/I0vZk7IWvcukExGrRxu/RgusyMrSrrAkyabfdiVy2kljVpNWveXnE/yY5/Czz5TTcfh8
TKiNWR6QFGkpPI5p2cnJAzXciehTYG8oY4UbfVGFgIUiXlY9gHDyzmC8sHQHXJZ0OzDis+uRLLa6
VPIY7+ZvP7jt2HG/NuCQhiFn98pserWsMAH/ijp17lgobjZpwvlVjWJjhSa9iD8ixn+K/ha1Btma
kNflj35JBZj5NO8Jn2IsDFtZ9fuF6jRhtsH1CjZ1LTFzTyV2ZXw225E+9VATuivwE0/uunQyaE1S
/EAj9ojiJ8P1A6leIkwSXtjtqq4yunYFscjq4sIVA+YdgKqjUwUJ7VKiMKo6KA9zDuOS6ELqCTMx
0pkxyCPbmlNFVo2XirgZx6UJWWqZFj1ELeXayRYaeD/fnHj/cxkO/aGbR66MOeHzz4p6ct98PCGj
Y/d/HIk7/N6hRjRiiYCpLdjUHhtI47I+uIQXupBk3sxPZCutVl8ns916qS5mFfJcV07v8Ixh81U4
mzWn5leYhXjoNgJ8q2RohL3CYxsVak+/kd2vptFs5KmSi7OjzOVPm+iHOy6dibHrB9PJVN4ZvXWT
qqprVdigMQDuxCYqnx4xkTOHSjDNB6/mPkDhuUxLyCmbD/uoPQCTlhHy/wxbVIMvRa+oB9qr2F9h
SHB458N8lh3JmPFTo3x/c4zHm7sv1n0Gg13xvZOrLZkNMKvP7E1BbnIR11FmbVxJ8QmuxvYxhw7G
qTC26vOHKLKR4lcBwIoSHH3gi5tiNcrDrXWZlkU2ciUwSWDnKk3uxpnF7BUUvQYrVPtTYgf2aF+j
2iceRHd0LsjaQo2WVOTsK9L9zGJKactF4Pwmn6pflyvScPItUDcHluIuggzbK1/RjzwP0KpBzdQF
V/IYWIaIdwqMnjMQs3jjbR4UIdsFBT30eE74gZAHb/mI73d0UAJ5zb9Pf6HjDNnLkJa0zdeLHyjd
wqe7/LjNUW4bdt9jVyPptrG1v9Xlt8aC9nm4iN6r3HBH6zxTNaazMQ/QYn1jnWovztIf7TGULtRR
SiAFjWObq+55xDtTATSxTYA/FQG+E2F3ocAXN28aAeTT6XtbLRaklZp35lBKY7eTdsZakJHGN6se
TbNVVdXMbNDrQNCEN9gOW40mqHluewdLVFhSNIQIMRru+sY8IKlK1oRQe4502of5Tl26b+wxmhvi
7Zjt5samt4KW1l1CuY/+DdsXmv11aAQ8OQPcU1HPktZQtr5LiDezlur+DX83sQdq+Dn+xDmTGYro
lFSAkk9/Po1HfEoOMv1iGC3aeFimO6Q2/Np3STUUJwG9dqYK7ISb5B29RmMsztzsaIxWL4OOe1WM
b1eBrVKMuUR7Y29Cvh7OaeebtNzrzABGQDqcsXsOH/YiI+FkD3sViUK2dVxft/2QPzJpsF2RGQLS
ac8bLfytDR2w1Y+M4frQF3BJeCAdy7vl7VsQXjM/lkqXJkZdFZsW/LmTZEFymkDieksQ1TKXPi3H
LsttB/GX+t/WNCO7X8y5Mk+8vSDN6eyWD8cY50g2VqLs74as7ZUvtbMnesG253bM0VAJEx1/+R3g
dRzfK6cxASEApOYSbsV3SpIuZcrJXpcY5tN6oI3biLymjy9hya4kLvmHRCasflQDxMhm7Yp9eUAJ
ER7HfdESUkFT8PiNY1Eoh3GvrfXabrEJE4b0jIchHqU7rj6Fuu9gForNZCLyThT/gqVw4pFc4JkM
WwB8KcodZdq4cOQ0S+C+G8b5M2Y7m886wSNMxqxT4OYDn4bOYe3d4qTBH3He35TNeEeWzovPRFjF
GImhEkHqNg7gEHiphVn5wmb50hQwOvX3IeLPSd7km33fVRA34ruko0gBtZGVijo+n2SDJ/oZL+n2
V+ri4+bYjqjCCRflGJz+fKXexdSckWw3lXUe6WzlmqdhOwDmfzwFGlgpsAstotLs2lAr5x45ip7D
wqvtOo4K4BKhVn8D2YMclTHc4mIEgs9qhp1i3nPd5uK3yFlr8IGT1iLokeqSxxMH7Hyq9JaYqjHl
bT8sbU7HEnSqWCYLfC6/EDweA0Gf/BAAw56bTqhSEzhOLpjDOpndTMzq1x8FGnhBjltx5zTQa4nw
egoJOalRK/KvYAhLg0iwUBMN6+QA8mL+GkwajxMUL2Ej8nJzVC+arIHREBe//ht6KzCGLbX5EYDP
YlG4m96mVQ1kiKjalpmPDAbx3CcC2tbnnFi7RWCUKPGRKwImH8Vp8AdU/cBVygJFRpNUUXpAtxq5
5gGzD7umdopfBTmUwf7JkbppoxrT8JD7ry2t7jeOYfc7HK9cSPztlZvnWd5AwZLejzdoUtdPKARS
zREKkJzQ97nI6sTjQwWcuJoAJpdW9ev1WhB1oROSg7Ke7Ecazb+39BrYNQ45Qu2nkrGaJV8W6VHF
FSnna1KKB3k6JyqKAV9MuelupWiNvQhT6LWLZNpZu3adrHxZYd5/z8+bZORbWNLKNHsKw64Jlk/2
6tjXchlxYC0D/XahHCn3BXlbC+/Iyo3Tgi1GYuIWGKCAsGWIsyHO0AFahJEgmJn3F/Tma6Kj5Bi/
Ibfxa8SdbZ8i4JW3nBDBZ6j4ytYv4PTcpfuDM6tN6mS9ViYaZTPn4PTJ1+GNcVK0OlYbVhf7BJ2M
EGopL793KxegfUVleNoQAG9KrtD8tRB0vL1+hKtWIak7stuKYG6LNCBhgW13AEk2J3BaogR6noKT
63Tak6W4bc8iTpcqky28PKGe0c4LGE9MF9X4zhq2Afev4yP/laGu5LsEdNUvwXcw4mzWJDFKYlu6
F8wQfghnhesy1AxSpwAzwydrbyN7/cFDfbW0dBSZ/eTIoGvnyVik9h49N3XM1SW2qKMOuODgFbbI
ibbg2LS5tGYStN9IY92qHiX5yKHH3TvT2nHtW2aKoZUDIoE2pIFd7MOgQ6/kNAN3KIDsWBoqgn9b
Y1VP72F4qOOUwzpuOEbNxn/+zoiejJzUMsCGneLVAEl+f50rztRfQJKuRHBI8dP1rZZFRP6VDdme
jSccK4UU/QTziPIPm+DRdu5OsjIcDmmSVaK2FT8a5juhdTrJPW+5jMd6MeFk0GkqpiODEixGPf0G
tPwrnoV1Rl27hudu7IVlurwU9SA9aOegqSedt5C8OQ4x+UoYxbcnQUa/hPsyCmo+MsGvPPHGoJ24
iBXJwAzuY75lPUxLy02piDsHEHfEma3vE/sldujkFDRI+XuCvN7qbFedhhGj3fAvYy1bRyUyhZnO
iqccuY60fhaMz/8ZF1PIBawPHWzrxbFk7s0XS7i+BiSaBogmQG/ZyPbWEnC0Mu163MfQI5UZNdXe
MXNDib2QwI84ZoZ/NFWgHYpg/PdSo2IMUdY+/CoezLx6qJeGZQuXrnOkn1kAKouZkJa34JJJIidC
Uzkkc5suNHBzwh8Sk8/+rp8zs/fpIjwd4/jbekLAqbWsuONYjxHmaBwNUXkl6vUh78C7mdYXLRqO
jUn8jlOpgVQy31Kx+yBc97+DHjsFVgbun83bbrO0kQ5Ti2jzH/CP6bckg7xpAwlQ0tNQeXeRxcla
Ml27sklaMsZFUqoBEWvsjr4zuK2qqqfTymsYIoTiQYjwH1vit1WZK/PhLQBuhiuiFQIFZ7lEfyvx
e6kCVNilDibwE2Oc4J2fOKv4vRcdR5yMVAg/p6u+8A+8DYYIN96aotPCH7zGCw/zPF+hkia3ukGB
U61AfYvpv19r+7+Uu/2EGY3oU3rPoC9APUw9G59+EWxj45KFszAqQKnAf7HsnMopNroWmBYzSctX
k9W7l/0GWkvSXC7U2+7lOpmaH4tG5GcyiGZwaQ8ustokhrhu9vwJMfpoBp7vufffT30FwleO5t0u
ifu/mLAcTZgjiIuGD2+hG85k/UZ5DHseFS4hI92f/oOzjbFTiItqQ9yOkUyjZf8aHV+SIApkzNeW
jxPw+vkXat7drn3LHhvWbqybKLCXkAAYVC3O2nexONSL+CgZgm7DxwBzQalybCrZ8H6Z0zGPngFt
p97/L9M683f4Sf9nyIGk6WtzwqmpPvKQzI29q5Iz5/k2Kt2csTU9Pptopx/qfhP5rZ6+bh3cwmdL
aga2Edr3GVxMdkybLMcuFvxh76p703cHvb4wJF3jy+5HOWTkapnC5oPDj38Qm2JIxShsfisvWGfX
UItM6pKVdEOjzzz/ts6McwweqDnmkBoiKLIIoOwsdl4WN5qboDXeyIwHJIHdg1fLj644PBs8Tq2Q
j9aHjeaEtAmwdCxuOTj8QXORj+6blrobKPz9T+LXvhEpIhFe/IR78Ii0GIgRCP6r+UHUn3GCJJRA
s2E4Ip7rDCuK0cvktzjKq06j8W2MtHet7SPDikNUPa77622AkzH7OSgmLDL9XPqW9G8gotAmtS54
6EzpZiTJdQKcSzcFYPcquTIRd0HonKcI3P7MTV8MtUSHMVA6Z/Fjbs8LlGEtt+1gzkxULC4YgtuJ
zHKwh5TkcSfQ0ZaE1YzHSRarTQX3Nw9oYikET5c/OzlfH7i/SPL6VhWStz0vGDO1C+WODgTNbUTh
h5pOg4wKHkiMrvusboBrRmw0fju+fYgoXr5U1WeKk85ofrVTGJCr5wG6fSyu0OtttS/Q8U18ZCtc
1ffXgiCb4c9ffQ9uZIoMNVDX8aHWmN85e8UpQ7Wfon8OGmc8tr5aYm0ggU+RREclWVyTqoDFnTVN
qgpNLhFZRTaJ65BLbNvawvpQCQCnJSStRxKkF/ohFn7IpIqs/oRQ9Jp65FaKQXZxEBQzUnay4KPq
85zGw7Ud0c5yh3thJbVe1Qv+XedSeKOXL0G+2WcQRGcIfjamInXKiWVmtFxcCREISQ7GhvFJ21AE
Iu0vIwgadWqDYlRl/WnFW+9+vVFbX6LXs6U8wSDDs1Wc59P1BgHcbWlaojHPLZes4mDMoplA482k
4Wp7cUuC1gMbL8mvD2DGT/L+YDpdzvs6uXpWak9FIvUYDeqozCeG7xhjFEXsZWQ7q3mmOXBLa1kG
K+hnyFwpVxRHXjKn7i2v+OvC1GKjikuFcfcZ9JvOokMVML08DZ26To5VWTZRB9jYVso3EQlWXBEO
cdSs9mFv1cFHXd72mDUvgQtdkGMhU5YyawYwPhXb4vto/lGo3lH1r2cIm5pa2eDvesMMRZVrfrjq
9bBm6k1eG4lhZcLWOTCUavi1KGDTk0fKXZCb1a2l/67xZAep56SFeJpQEt7kYpfeYGlxpU0TtPbR
VdIws/qX0ISCzz0BFHbs2eJB0MeGiRms1/F3tC4+3SPkk+qyX8Ut7ajLyaMsd5fsSowJGtLav+Pd
llTYWspY9iVXPblRX+mB/dXcBQAcUhwXSo2TsU5LAfhRYIkCy+vkl60CBy6nfoi82NVFL+/Uh3GL
xrBD/PexT8+kTCsJ97v7jpwDg7SQ/Hd7QpBnCtfOPWWRYTfcOHtUYp7ve4cCKJCxFzlfuFqDbAhM
tA3VOTcAGODhv15xMmHlWkZx38LuxJm+mYXECbuPMFZF/GrtC84kYc+tz/39MyR3p0VZPOTjBfDC
hetwttK7791i3k+YR+YOfvwMyTqCgodEJbi+dUO8grR1TPUiWgcZSmSLMtRwIBuqw8aPu/0nL0rh
Omixp4gl5fCyOsVf0O+Rh/BZ73LY6AlZtOBzH3eZDfy74P+MxVBsmBCXBn4mOcJzsGc4ircDJaQl
W9zq34geLWnxH5RZy/XNJ/QeXf0E4OrShdfPgvPSDCA5gbWELcX9lMgpOA3am63GjBDJeSpsnEwv
Zxtts/KW3sRMeej25Fyc3Zh+PrR5pLyHi4z8uVyoFUiAzWr1x3Wx8G8nClrynNzxrjym8YW+reCy
tBdoxeJfF+bbBuh6QGdH/7LVfhDEGnVEjv0n3LFt5je5lfOZeZsIZS/FT/5lNg0DnIJj3zjnSZAD
RZDd+bEodHHmZpSM6/Bau6SsA3IXjwYRikewGHR9coy/ni/tepAMibbNDwSbni8A/OV1XvnybjZp
Wqusy+YdvRcJvGLANMhcLMuJbNWPx9ZmE3R5ssZe7K7y4EwVGQkNOfOIjWHthQFG0im0OGXva4I/
keB2tnbgibstaWSmQERb6I0fJC5cHTJcvTmCsAmpnKGOue/yZuXVQSeowA1lvyuDTSerwwHupN/X
ztPXovpbXU27IQziE90IC3hI+gAEsO7TVF3G6lFdrPyKX+92OLkKqDGuOhPXbsid1qHDFRNRbYNv
LnTC3sVMc/dk09jlD5UJEBpAJmQrrc8HBzCOXuPGFmfvHeE4D92snUrabvjHwH/4kgy7B8OAXcoW
Wz7BuriUNWhY14Klfgo3Nqk40O5ELOC2feLuUdagz/jyxAAz84lo9f82PSw1KHzSXvxPbjireZat
61HvbFtzlj5zS5p4mV+Ispz6Yo+pxRkWkc7eiNt0L6bNAwBba1veCSWDkgnbcMKlv7DIG1XlqKL3
BQgkfidx3t92zIokFqkooDY1RWD0wv7tW1VBGni4+yZARXe9BM/LYHlhWPxZar/r8XViwKPztL+u
g7vTdD/YS4kfg+QkyefcYjXM7U9G5Xad4w/haoN5Ideq7Gaz7OFn+YMyhTSxOPBNbbnF/ragzGi2
GvpIztA631ZaNktfQO41aWrlCvdwqKdfaLE+i4ZDvOjtnY2W6FoT7fsibBZ+8ucCSAVCpPOoI6jG
ZFI2+B0FUaexIzT0svsxtn+F5kkBYfPckyeQvaAMLon+gCUyoXYkM6lU2lERAGFB1/PFSmZW6U0f
Ef6a103XUfmoSKbYSRHOZuPJyg+onf1y+EO0S5rg8Hs8E+XkEuwgBCU2M2UAZUzazxWXUuq3hsxc
ecKYnK+/TjpyuZFKqCE0WCrCr4IVTohNgi8ZM7xWaVxf6xgcaT/i6XxLsOTmmWLEi67QkDYYh3s8
yHG2FGGqDTAyEUfGaf5oiEMMChpbAuOmcH1eMtKjuNF+6xwX2gBIH2iomGnyVg5VopMitwik7KWF
1nWkEGuqWxDAtjZC7nkjmPiSCmi7OvCrt7YXmIFUvyfcv8fO/KGFAcpcz40rtzVFzxi1RgY5ihwe
d5MAaG4LzEHDmREFjW/+aDJIH7unvTjR9I65WZHysEFSvZ0oBbds7wHpxq4FHzqjh9hjWpnp5DPz
kjw7f6M/TVq0M8zlURfHPcjZZr9w9P00r2bBQeAovmi8z4sXkLlFda8DJ4PRa3Y1AyuD2mwGMq29
1B+VgELwIQ5HFur8dbI3SvovG1dfQzRy6wWyM9MUvfGWHZaOUswF0BS01pPWzZXkw8yNvQu6rlm5
nsW6brNryf6UtbIZK8WZvnlY4Cmg/vR1TYgBL7V5hPGNR91jHl9d3tbatrRgupP4k1cc+3t7JfoC
6gHsQxj8pMjqtoPJITdZoT9YWhfyAl6Oa10MrDjDSC5WqWPax0qQPgIjANBlvaIloS1BicTfquUT
lIWeLjyi3kWl1EhX6/HWbmncmb6Xm5gkXUI2BUGvQlBN70Er1uNqRFVNP0VRdyME3YVSdxRZ0U4a
fn+BLIY8dWywm9+XqVfBkktgwrm0fdaJNvhRM+OlBTM5BG0Z+Uqei8Xk86/Uy1XTw0d+VTYvDAYf
gQIZPXlzFg3Rnx5B/hFvv20JvR2W80RcjDDIbptluBmw2TJmvNREK2pHOSJ7RxZ01OUHPt0hx7C8
HyHZtDF7VMWLMiRnEQPv4waRlZpNMBf0g+BedY3uNKTAetSuxO7H8SrhH89KpWrBsFa8otrE4LLe
8EYiTTb1MH7ggDXTIq0UQJDMTuOmaUGFZVspCqVhgaU1L1GJ2gyGFkcLivgxR9LZM38vebOwdFXI
60zaoO0M4nOTdfaFvXKdA0Lr2Lyn4HSpzmx2gf7AtJjlshf3grJkNUSmNUnZOTL4T1uTnrKYnO3F
b3+myQpVORLx5E6g7KMUpjuZUPvYMYUN2C4U8N7gF0zJYE6hcofRZ3zWEf39AtZxpCCySrcg7NeB
uCm8s87fnOHvEFi3ihhI/hJLbenxJeV4/mOeSKIb5fGEpItNmO4B08AnNVCojsJunYZLlkks4E0K
pqKd0gHHCDFbR3Rc0Hnm7HOw1qJaP8SMbKtXdSTL24gZc/s6NIv7oRME4bsXtSsJUp8QJzXbU5gN
AoxnGDKbaNPtp4nQySbo4dHfm5a0ZTFmbqaTTLmFaMDSZfVPmVB1dfzkTzeDjdz6T/KRV0vuArf6
oqG1rQzoLd+jSX2x2KJOvZ8soIkg86Rl6Ds5jaAWy3NnIjINjAaz7Vk9eqg8j4Yw7LAcL+Pm/OxH
6iCzieEK3wZOwXc/pXCOWByWl4ZOW9ArlwoT/6CfxgxL64FMnvKP+oJ8R471XehgyHdNyqh1AGEH
guiHBpHz6lXtZd0JoJXNUBHJhCrp8VTjYpR8p8QPlGnLKl2lzoObBO6vU5ohJ2ePyWlNwLspm/dA
zsJvjwtKzXeSgqDaBo7Y8UqJnrYoEepz61rZ6Gsb0bc5RjXiYCP51cBqgLOFfpUbB9vyn7yJQy/p
K3ZhPRYARPO2q19WdjHZcCLmBEBelgIneTjazm1CAv3x/YQfb8J6M8Qyrlv6PaOkCi6ZDFefLK0A
moMg1hGrNWfcZQOvQYZk3qxhOtZytxeaqRmCUe40cEUssn04vFQiHZvJ4CLVrmveG5GkR5kZy0YB
Gpatv+84MDydhIUHyVZ7/vYOnfOXBKbbS2PSX0Emu3da277rS0LOkFSiWxPzEIMdovUuLhpYVV4s
+ILfproDjwP7+NRZPbMctBiKPteSRWp9x9ltJVOfJG+DAmWo75Ucsv7yV6GGUHqptSTp9Yj+pPAK
J3pwdYQWim3Lbtqo8BKReaoLI2cqHlqzOOkewkys/ttmx+zG1NM2ooTDStfxD8Gmr2XZjJevF5wS
KOac2NY1vaJF1Cv3MNgDvum897TZHKYRICO3efZlk7FaM5Gac0lR4tA+c1VetwMRf8HAJzK+Daba
0L++zr9ZzXtVNkzD3+POCf6PYWmGqW0Cn73j1aUkf3IhhrY6LclNu7cKDJGOf9q+FtMbGedfehw4
GvVY5CLALifsp8Q/81SCn9MHPYo4Jl2CcqHVtZq+IUe+k1e23udm8rsX7dLNlkkmsz0lXRea1K/0
4VQkK/a5Avu/yprWIOSCw1kX4jtKPvY9durm5y7b+KTSL7cVz0rHJw0yEyZSUbLBg2iQBvdEZ8lH
/vgCZRQVgtE3jTg0p0woE2Ahs0btO/A+wkOSYYIAy6ZdfuJJwf3075JWBYYfMnNJItAdDWuxEvWx
7iVzjhEzd1a81MvABCvKTnjL5F2LABYzQqNwWSOcUR+Xr5EIbLQdbdDnhd70s8MtzlxVTIjuIcWU
jZ/R6kWQvpnPkece1rAhkQWYTbiHYfHLF63H+obzRZO9zDtZw17+EcJal/qo7mWz4uYpECtB8HeM
HDxR4nPcJHnYqWNliTGjZ9cNpKrTz3nEaTPEaJ70+5OVO3bYBjelsCKZJXdAZpyHbNGwAaQj5EP7
W5oiSFEy2ydHDnXP5EOXf/bf45OpCQCnnq01WoMeAEpbhEVB0t7C/zfo6/j8RCdoCYJje3Wg7KxA
tKnMqKPPzdEhxzkdhxX4IkA+z66vZ6L70HKPBJyvwQ9AJonuoWID1GtaighkYHeoFN3ThqHOSkSU
V6pNAO8QluAT5AFcdsblPCGkEliGZ1UNmq2zRpJgAFKGZz2NIgQyizCpilsWL39vDLwk1mw2eL1n
ehGAEKpWKQ/qWlUt9mK0E0Xy88koPwT6wc38UJbFWVHUBAQNgml5VdyHbc2vcicCrQlh4ITlnQGc
BXS9Ooako//jHnr31WroJRVoRnEM6tPnvSh15zPrlasbFAiUTJ6ECpFB/R3V0VrBwFghGceAgLLu
wVbCFhIK1fXzTOFMgsHIxTV/VnOztyPI2rlAjzsRBgB0La3TicSspyo9wx+MD7kwJ+4TR8gZ9MD3
OQecnGmHoEDa4qKX6A7HAMYDXa68VI+TetbHrYzRVENkxpscNqPHVvj+iVC8rR3sWmaAYx8BjEdV
FEp6bpPkxhll9CtilfuPY/6WYfJjbo7vT+GUGQrOuLVzERAt5cwmbL7y9meVjxf+9S0wk0ry0r8Y
91rscfsWbRjm0kXmX4Q+B8KgB8dY2PqUoDOHpjWmmIKK0h3y90FSstdWlWlAX3/cJIthJLca5EoE
8oeW2x6OAtWhMC2ssKExmGxSHqMwZZl+C3EwtSNS2sXkwq7yavRwhuSTw3TSqxtbt6NpwXrQXiGV
hZkoJxR76yYsn0DMzjhJJ6sH2vpwexA+62wKCNPvZccFzlsEeAv9KOFzeykMfH2a+nx9kDVqSY8g
btQ50qkg/0f6T036mEab+uUjz2ciS0CgAwseMlo1gOU7WBHHJJ8MpHBtat7DOkRxIZkF4YBd/HSb
7iiay6mwdl2sAysvnEVg6CH3If6nEqdXIjudt/2Fi3Y1pyH0TXk2wAe3eOoVikAjq8suc7SYmYbp
HGev1wM4qq8/ycnM66hh3w6TirUWXbNM2WBn6jwOORjyjCVEmJky796mna1DVb5keCdWv+1FEx21
4T17yPdcNe11ZmLiIHp0ixdLYpDyM6Di5v4ZcxEGQKFadgpzmeqh80HK7/K70j79MsNKckLYdSe4
RyHhcuC4+tvNCVPNGTS57TKkqSdbT3F3AFIPv/6xBFl6Dsg9p9LBVonxSgJq40zaUKFrJQBK8y3T
eapIcoMIoNMZuXqtBGHx+hVH1G3ZK/528bA08Yo6Ma/9NVGf0DM0z4E+Jy5bBb+k0Weexx5WCB/l
cZKbm8s4/QgAXgReeDy7Eg0PfIUJZEDypI4vbLmK70ILH9vvQqQp8zkZ3g1+7Fg1INjtg+XPSWSG
ianO0cgoply83ddZtcgbS9sXDZSfEyWjr0DD6H/icMel8S/bUb8nZ9J5W7lvi6nbZhWFeiZAJpbW
kzqySlmxZMvePaZiWMo5q4EIN2j3jAfAnhmeoBhoK/6hHPN7RkA+zE3M9pJrGBuhNquDUpWdL6jN
KxCn5md343k9k+YFSrt47igLVanrosR4rFgi83ZRugt7eybhgMyCZeeRyEauum4sJR8uVdUEME80
e/9Y4mVjUWAB9guxbgTFIfX+WDT6zAxqhkuTyPCZ3jkGwwph+lrU0Ebu/v42CPNvpnOsZW4PcsMd
QCBP77PTKMtgho0cocwTHxFO48u055R5pcT3ISymlv5O9+DyFMTtdQL9L8kq68tSifaHGrVT0jsO
0ZsHe9aKgTaqVCPuc4QAMAM933o5/v4q9aqzItU5hKqHQafqO+4I+fN+skFK/hzdiWZ/bBMDlvaq
yHgnOBDTh8+jPQV618driWrV7eAx60Ro14QDDpn8Fu0eCeWdwSXYOIklcyJJ4aLMCS5ZFEqDi1tz
V3ODGcTmgCYyhRNsmWypm//RDDTV/W3SIwOp3Y0i0qbmA3UGCjtC2Dzy/n9cA+t47WhWtFyWZCwN
Ndl079X3SFycQOcXmkMVTo5qZvrbPDX9M1zcJbLVnlMsvMP1p3MY2/dmyk1/JIovHwJGZ5dh4ESc
JH2fS1TRPbFP5zDCdIl/FWDeidAcoP2sJ8ZeZFYMFTCN0KkK9XyUwzbsldQYDzfeOtx7V0Al5wvx
QTAMj1XiaiI3pLPS6B4vKkLLlB31t7f4YrRMKMI+L7U8sl9fYe8DM2j0gv5n3MLzxhQFkKxC48UR
bKXSh8vQBTlv7/nbxvio6SB8YPXm6tizysfoThwyxbfqHX1VLX+3UBqCXph6djMCF5QnpEqFRk/V
ABxMVn/TliFGicYZRhWnye4kySBauyZMDVEFLZysOj4b5W9ZZcg2Zpb9qxOpQxzKHxGZZczDLg/5
m4/nMAstEz1yJMFP7aY1Jh3dKaUjRG9exkRew/njH1ct5SEUK5WU1Pb074eXWSL5MVcwyGtUtJzy
a1FlADJbylsZJpYn98iYzhySo7TUOuTIVG7Ef/pxm9XMGy1F+Vm6idN3FUo/r9mU4un5SOEouYX0
X2aUg6JmRZHL72wB/sabqdKXYVFgtsX3GN/kCVhWD6+5qYRb2HlaorRdXEcABiiyCrCkIZnVGlX0
RFffv+9Cu27nH6ApUwp1PDzRHOSGTBIfGuzrNRbjSNfpOfenelD0Nizb6laqZ8ZoSoIwyACJ8Grd
0HJaQRgP4Ls94EgKapj8UK4ev0AwYlvOih7pR8OFLJuosEXE4CBE/JhKJRzhqLqhfPuedkxxH1bL
aMcf+64MxQbZkQtl2GC03ivusoOYfJ5Aedwl6l3JVLn7LAP7Rpz/hUf6tlTkTREwp7N2uQkvfpqi
KW0wpHCuOhLInzT4FvhAeTCRhcEM2RKMBrAzCaz1rZQrebPIVybYAigzANonL+kAWz3MuwWVv2ZU
X6MYcQCsJvrzfmuuADWVfn1CE36E7LbX8Vw8HCdKtDNur+gRn+ZUoTmHWO5S4ZdojUINo0gDRi5O
t8hfiZldHckDuuoS/JTIPVJfgxxTVl38cABwtzSeRBIHZ7FN3V5Z6eX6WtPwOU7KXuPHGoMdS9Yf
9MYFeAp0y35NH4J4dVZ7J95nWcwhdXW9JbT5xoV2ayw3Wb56ZYa8arl68zgUyiO3yVsdTmitu7u8
tsOQQIKTAVbM+ocKn/QnB95MwNcUfifl0kkyjwbqesc6iirGxRPT/CfWTexUClxW3ORvWVzlonD0
ce38n/2pS4yj+mEalAY5EsEicTUnf5hoX2/mOQB2TrGOaYqNjoi+t2nAfEyyyQYTLCyzHHG6Rxvy
E+4V2JPfXkysdrtqc8tUL4ltLyhYxpAJmj/MiCpafQRGGWOeNxwPgNxlxSM7D6/6OVouwpnqiQ2O
m1OAFCzWaKSVym7mX3o3FpW7jxKajQ/UbkJvtgkeRRFaPGh4YEY+mJR7ihtKlrJ1K5F7OX+li2hy
2aw2cgZRUKjb8HbkH/ZKMefDk36saE8Vm7T8sLvkleheT0BRZ/MFGyYrKKB2hjhQlWYkwO5yTkok
6VrsXZE2864UMH6pFVa3Kxl+d7kwm55u19P6gRfwhcSm8X8bBsEChZIiaHyRAQ7eG38CsXsmGDD5
R8njQYY9nvnjGuL0Ics1Sn9K8u1dVM3UQr5jk2OTZ575Vsf643+k4hGNcQ+gt4MAWykHzoIoHPh2
5S7xxUAj6WSoymElnSPkPDdoS6t4rxZ5Xoc1vVH4d1g1+B6lqtejDxyqw4LppbpgqyIPoJtn76M2
7Ft26Qm/iixPY51ma3zZjmeuytVV6xMywNZA0Pz5dqadpHBgDXYRNYJnJbDoDD+ReLKf3VskbIlb
8FWQkjuSTpK5B69RY2CTOk3CJ0RsB9nsNK72VkZgMCy+iK64CJzpf/VSxw3HJvVMn94porBDfb3R
/gwY0b34DYP7KvQKgF0OAuUz86TL5ORwC1A3u/AFY92AycdFhMpZ84JGjq9bMzuXC9srdaa1QbMJ
IIGOKhxfMu1P032eWbD157o/6pEgyoLCq9EE5bj1uFrejDYFPf05DkZtOaoX7P3qXR+753IyPk/6
iL+16DX81OiIBFQn+RlwT09gysC4xJKLAbRpxduaalkM9E1NTs9eQ8TDxNXIi8GYr3K9wah7JJif
XioZT/59mkyQx0mpZKu7ciW+1jDWhaJ7yLpAE91hF4x19YgTlWjPQM+ekSQMlil2lskg+sa6JanY
DlWD5G4tVQ6p2YSyWJwGnuY30zJn7FGy/ZUTRE+rBWH4D9+1EJ+Ed8CPGFRe0/F1oWW2Axp7Gx3m
vAzgxGg+7Wr7R1uwVbL0W28rg8q13TuAzbMncep+KNMWP/6axTnMqi060pAUWVQL4N6Lmt2V16r2
/IN13vun0YbaI52rKeOuOf+r1mchJuAdlwAcJ4SiCRs7OQsJdBRRHpPepR7j3z9UAQXoXTpindeM
NBjDL13dA4ix9u2MMTrqgIAeTlz7kIANK/XjDUIxm/MqhGCpfP4036lZ53uVxvVZGGu1C8oZLGhE
Vnbu4eVCf6Ti8r/24/DnCAS4nssGUVYQUHCVq12XZJLnINTdWhxpbvkyBeBwkiZdVdh1IAwzlEqH
z1EhhoogWXvvWUT7+8rPMtaqGv5aXouQQLafVGKgsBaqa65irDBI8SFJeVzHTaej5ETz10fRdyzV
hws1ttKkdDzcjTcn98b6cVDmF9fDbLm6olUNXk4srvuZ2apnHdGNmRSWQF9sr6fnlENHXCBXGnrs
oHSlPp3C6yZeAuG7WCj5Xnqpa02Rs271uTaDPwOdrgZSnn9gWZo8A/fCYHZ6uKF3kUfWNXTLmdnt
y1Rvb6/V2GLqURiePUsmJcF9Ldm+A80lLfcPy2cUAiXcqxIJ1bxURlxpz3DTB3r2oKyegOzUmaOl
xlN4+2MG1f2If6vMx+bT6w39yZrFa1fs2EB5fs89tzhFvjdU5ZT/HabAJG5k3dhpchzSpgAIT/cU
kUne3lva1grUYO15X17adma+bTvrE08bX2CzGgqhPtAWKvh88JTwrhpfpdOPYLFvEVANt+nfoc/z
QiHfmBzojUi7SPMkw/bjaKOeRbe034bkzZckcaPxdx4/plM/3axlST3wKKna2xZ+sI3isS3qeJV1
dPf+POunr6t0ACEmVIiF0d6DuRLSiBGueTBIzVGMFTU1lcEqVZ9VPBrulhvKJDLgHI34kDFmDsV0
n9z4V0EFpXK9bJTp4L+gvA5oV/pLKSP4UWJ0zDeCNsI4d3hq5tLSNcT2Y+QMH7+/yfOyBjlvDYXs
sIcdukTwMxyvMZIwV/ffmzzE2Czaauurlk8MY4uj4CMEb3G7HTFFjmszSTUVjK+eMRs4ajWb9/7i
K29eo88vxjHE72/xMGOUyyRc/HgEKpF2Jz+4xlq71gWU7kl6mqSj5OqrnF8ZR86BqrJleQRKCCXM
dsKoWx82YGnpotPEEsD4Z4BysJE/oP1VbdvBQCGnwz5PXfbZnkuHtiNsUt6mdNSXGwQz15tvIYDD
zy3n++Y3CdwxyL8V6BqV3BLDRT0sdjWFtkmkByMBw3o7Qa0b8y2UgfGkH9xBUqTpDBEgBO4uWsW8
Moydcz+2132smDKFCQMqbnUmNXsfLmnOpG6hVjYJESPqh9/5F4cX39qy/bmrSimR6fALzCqN1BDi
BA7mQKKFZ5PODd3BQ8KwqyHs9pvdyV/7d0RUprStcN15IiuqesfmK5ZfhVvEmXJblG5LHktzLDuW
G2kPnhAR/WJKQ3E2ibBeChJfKnNYjS4cj7Alx1DPj/+9WQT383hzzc8QSYcy+vf2Cf8lCYHW/7p6
L+AX8TnJ6H6qwNmYEp00OorFPry8iXbomVdjUpXDcuTz26iuesHAnO7tFV6ZRihARFiPFWu6g3iV
inZoxZysnuIA3xhLBS/JYiejlQuoWUA6KPND1f/epqAllmyGs1bIgNo9cCoPVwDjmZIKFwcS7zh7
n0Rgn2rNp6dpzIssXgB60L3LFgQlYoGyXa+Gswm/LiIbuU18EJNLcylkMmwWO2vm3ioZ1SR/z0zq
wwK1Y7e3TBy0bSSTwiVncZP5IjVR4GPoLAEImH8D3HCZTxH8Mw9YjcswFDh7/9vZIKihj3E7r7wK
A30zRIuvKX9YyaZs33uwgxvOfdt/9s0rLYc3AxFmR13EZVNMl6ox1fDRLjaHwBoI1wGQ4tv4uvkg
zRaZqZAuDUzkYQTwcHp3Yx/usmipRIAKKE9GPHUSABknUigaRLYDlo3zefp3maTtgspWyboX8gxv
vuFnyySO54hYbfqGvtLWicR/SBT69P+kCsyQlQYN+W60zZAHO0kV04r8K+4Q/N36sJn8FE2xWtiA
jcCcg/TmwMPh7B+5T6i+2n/lc8oqS453q08yZFCB3m97i8fN9NoSb2TOIRXQgr72ZAesiIQSoLzS
6U1s/Tqq8A3qAlwH/4rVG6JBy8Z5P7kOtnPjbflUtb4BikuWKm52DWkeFj7Ap2zr203mcgztGcTu
hXdSbS+zbs76kzCVA3Nq6Id05g2p/PuxtSYFcYIbj0jTQMfB74JdI2cjvAhRHbvd2mFCUNlIdmmK
m8Dwpgj/LDb+owywsKEAg/brvVXNrquSw5kq+6rEZ9Lfp+VjirEF9dXrf27DKj4QiQTSwMn5MKyw
YYSBxThMKhRIyzUvhy/++HnxzQpzBuyQtU8LaQzUaKs7u27FBH5+RRCteXzlCMciobyksoBZzHw6
AYhbrk12fiOblLWthnE3W+BvKR5fc+beME2hAlwvpoNwrbt4mJsQEfHA3T4mJq4FLwH7lYV9n+0z
b8PvLLEyQoLcTHsgUHaOI+RXwyCCtAZ6wF1T20XGBngXOdMmct3m9lC/KQc2FWtpIINyjyGcKF4v
UoAtHEdHK8Pv8djWKZlnlXNwJgMZWRmdvg8ZJq1CvaTAg7lOckhuiHm/yL/d/jw5jL/Xhc2ygBOT
aD+zejD1et2unF5a12ZpO9p3nXWQEGNJNli21HiWhKinNrQy/1p0AIbXAZlR/7Nsu9M2uWQfTKuD
ElTFNF+hwLMtRCa6INZNIP5olVdQ7RyAmKjLsQL7PLAQ2V+Gie8D8wAget40tvOD6WQfcGgJqJO5
Y2V34Q3djRb/Vs3BeFOSUaMEdAPlxU+wdYOIgJFbUTQFTZFWWSDh2OYUio8e/LeRlZM0H4Ky8bKl
7GBFXznqjNVQfs92DOdQw2T2SHbpAdkP6heW+zJSpOUQWlvaMrbg+UqPdusNTp4MXFPwF7QtDdJg
oJ2bMdm1lfgewNZEYAxCQMoSnLhW53BpXJzQeJKwP/Z/fYYfd3MOYJTl+xQRHa2lQShzwXz2Wsec
h0uAgTosupMn3MZJqmJ32NQYZ8F0oSl8y3kSLKalGXitPCiy/Ju2CTThGZaj9v/GoD4FOZylz/do
JGNrpbd5D3KowBqQP5l9s2Eg96842xLlrUg6VFTDo8cVUylIoFLS/Cz99y792cE6rTAdbR2JzlTy
pZg3DpCrplZ3mVRw+zc2/IoLuGfr32Ks46S0h8TV7qxH4gtFOGzSwa8TrDFLB88/P0u9Og73mcjd
o7Z2iO+Si1AjShKHXNwwB+NLQsS32kd4VXOkRFXUBZDqtcNKQvrry+H16NaPVpD2uyAREo0rjUCh
pMnsEkE9zSHFb1CUtpf0NKrvlkvMHHb+QTNGnVn0RwyBAqs1aFSIYJNoEJxz5p4vpas8/uwnu1+9
MuI0MpR+oZI5NDYwuXJil2seEXhaI5wo2smDFkgrk8czsNX6jtv5NvFJ+RSU7x588g2sRf3BZ2Uj
chNqjHTKlIWvkeKylTYItTqFtC/EmiDoQ3Iohu+sdKIuZIQ2dyt0t3x5+2nLTLhUuRzAbnGiNX6D
ZRTg5Gt+7DwZ1jLnxXMrF9KH5Q1R0OxRUihxMgD/RND3fiXNUi80mwErATu/w8WNSNaYVkbn3LV1
gRPd3RWgQXdjy2Z0VmgLqBi4Q/JZZ0Opu6Jz9C7BBMv/zQfDAY0l40Q4rfukO/cwJ5TqEWGRbV1p
H6pCXO/UaxpMNmKsCUSUXB/d99Bbteqq0RudXmQfue1FyyTR9Iv0wAYw3RC5zvyGPKoNrbg0EuDF
wRrDjJl/dSOF/VfeRkMe4YnB8QKU5qpnalvFAmWAkVryberUqsvBb6mJnLQ8rmtprnGnv6SLEdnB
atMHPvtYXQwNIddTfPNo6RhHp2Fs07ZTbNqpwyCFFCKvwE5mcXmJXT/dBsaXgSct+YNgxr42Sydf
LBVUs7Vm/kLa1542B/jpWSR7uYSigPsN4uA4YbjAQoP1u8STrpIg4ppgZ0t3PGO9R+aFs2j0NOXM
Mh/tJnZHX0SkRtdtyofKYKFVEYg+6mrz7aav59bCLBJyq9OBOn4IZrqZjixIyDgRlX/6bKj4m30l
ba4O4152oXqEor0FbJONZrWmGt4YW3+04bJXDOdQgb0bgo98D7icSJF+3+NoisI8+hojUThzCAdr
TS33+e51L5wGYSlBvy2U0MomqSXQVze4xxKtecrr1FJY7Si8tVKr0CnDLOY/cdvZniKlNC9nC2cx
z+rqvYOLGsay/BtDbHPX9St47RbpCw9zl/Ag0bYJSGFWBOBPHf6VN/G5x5bYHr3P4c8u6GshHdcc
jQtvwaRuRCW5UYuNW8BAItn+wgPNkrgj3Z1HdykHr1GZEHmkLPRk8cF5MA9+Laz1gF9674eTWOa5
U1DZyoeLzNd8BxAkUliZ0CkKwR/syUnCChdqVh/KBbsIblsDgV6d2TS8mw0lV31x7AIn+rEZc0Jn
no+tzAbaf1QhGls0Yje3d5rJY3zoP29YydKJFx5sy9EIb2mSKBd1af1QGvW6nz9RG0GaOnIqMQ5/
JG6/WU6psc802oXRnmEh2DfOPFaZIBAAZTu6hzUQpX9oCouI3m3IpP4+8oYgXp0TwRcdP/fnk716
e8ddDqgOiMbPMw5Hgb4VigQ5mpNNJPFBWsGgsFD/HrBav8YwYL0LuQgXWTp1Z2djcO+CqixLK5qP
eqUJYSkp6+kHQ+T8JvUZBr9/4DQAC57cX1frXiLUcVsPOrzTBz7xdcsbQC2tZ8bSsaCwrB/sHCU8
BFcUN4+w/2ELH9B6AB7R3v73cQzt/dG0KFqyl6bwnxluvtdgihIwAQiM/XXssQ3ql1opm4l6TtPB
27VztH3lTX+cN0aB2aiHlSiz9fbZVCmOSzjkX5NyARsz7M7kVnMdyMk4Cg6XFHVICBnS2ox2MQBr
Uj6JMItQgMj2xR87dNF6DjsGcEkvMyBsvTby6Xtr5fU6W6Ggb96oSZMmEHv3RF4UjAZe5LyBShLI
Wo4hrrJfjS5trmsEN4uTtNyZdwvb7qyrE3e+9sNO3X/bb1SIfFzRzn7N3vM8TFP69LoF0s1IYlQ1
zs3nbCHaynD2ZyRzF0PcKWfPjoA89PObX/2+aEMAlnFG5tPDMt5msQTO5lGVBI7SaVATOaE2RABi
rXPqM85ZP8XZ43E/zRzNajlxESvTCL4U+qMAQ6QcwwXNLtLJitP2p+GC5RQ/Q8B8DIX1/G4qrCqR
AbzcQC8H+cJysiO+NTtgoGCgp4pU0KamaU36xC0uo9y4ly77Ge2KDbFXg3sOniHdQcU4Rgb/cUeg
D3b12mtJ0tX5my+UVlBPPWCwo04jvDBaVz4Tbs1qiSKoX9W5Y6iKa0RCW1v7THcjfMeSsh+zUPK6
Iur+73Znn2he3i34V+w08hGIWxGhYbyiIrq8iCaQaKKMTk2Vb0LNZr0kPEFySTMHxBa0q3LxQZRb
wM39fck59iKpGM16qPbHYQ4WDx0coTIf9aKfCc5/Wi6KwFiRHF/AJ0MFHKVqQBwjd1hQbNsegLJ6
xlLresiAXm31o0FWzQai14nR3SRfugIG7ZYeERkVx+11GOp9okVwCE/xWXk3y5WdZE/5DMsfSlYK
+LrnbtmQkwMEMxam5/JDXmEYbiJHWy3aDXFYO6RorpAz4radCnKbg/7dpWPy0tQ2KJZ0dsiMxAS9
7AVc9Fb86oQI6961U1bM0Qvv3YHZb4MnK8YCwqdxvXqdY5kt+h/R0YZpRSZMBiOay9pcrOI+rv+W
w8BZlp9Srqu5xDqSniHy8qCgvOi375OrXWlHsVSEn9HDFJ0GwdDh2RcFWqwl3Vy/a+Pto2DDwVkk
cNFcKKJsfbnsRRfGtNCacbS2uWhjfbLUtw43BK0eVc0+qhzu+CPvF46qJdDiNlGj9iLQQm79qWBj
rFY9JvMrZGDpV3ejwKvzX4cKARwfNJ9wwKbOyqJOFocMpC6QFYE2Ek+jEgEs88XilWVXD/f3NPxS
r6Wv3QVVnECGyAF9kAbeTex2ZzeDL9gM6XaPj86efuH7oE6nM56BbjmauAtO/NW8TapkzLMPaAz2
FA76bD7E/admq8tN6xZ22D7XU7dWM8EFDTpuY2327VvN2D3Sig/bK0D8Aw+gmumYhEHOrzWBO+Er
ri03f6KaWOOGf0IZBoQIYzLhOV0/gK+7LNL3f6aP9GgkqxSrasggPrIWaLUuWxaNFxvTQgbPX4d6
OQRmLGPmwJMI3TPXF6iKuyPNT7D7QH5iOI2veU9CdnEwcqXvkgnGN8YCsvOIi/naDRZIW0NrpSIf
Z0U/rkv1EKqcpPZbOqe51YxGHGCYwf3nkM3d9D4qnfU4Wb3fNboSS6no189Ypxqky1URJPR5E1rt
YfrBtMB6wAaaHzeb/jV1nCIYfUIaUXIutJQPt08n8TENUfAszQA7rl5suAtWM8r8uQ3AwsE/pmn2
gVjLOeojzZcn/lsFwnspTcYWDwpoCIWmCjoSYdC0bp+lwnsjmAEs6iAlRoQ63OKZhlqgtXwy4XcM
p2XV2beB1FAv/H6nbLQ7VdvYfsozt55jh5DcN86wgj5wp1Z2eEhvTjVC8zS0Rv0/FYJswfFbqnqx
0i1FjRnuPUR/c2CNst88kZueBLMklZWoDU5cafdr5NnBszdU0GYQ3YoHCw3p1SttZUK40IJhgKOM
CiMW/H2tr7j4sWN9EllGEzWZz7XYhtaCwzLfwWMIolhkDJhoOsaXcY8T9SKN6PUptZWGFSANd8JR
WYVPbQOGzeuLhivz1inioXtyjT5D64ntMhGcT/8u0VNrvRMalDCuBnsXlQbNKLmJH+3JIHoHMkUA
l1dm2ku47PY8CrawbecVYyu+HvTbEg45iayB7CnOmQoGiEwmUcDhGYxB0Jh2bz6gQ8F8/ZC+RAOy
RP4psBc1Xyk1beaPEPtFKBFcIQZ/2Big+JHANWS0WbpOomC8E6aiKRiieEcgg2HgbfoIfnXF/GRm
iqh38sOSPAETrVymcPFml4oi3wg77YaRWs8pjrATk2e3kxk0MrohWeEmgZcNX0evc2oFhKDL5vum
t6Y4o4sttp7Rk4BzuHJ4B6xJIzNzK5TxdNR4qPxWUTFzcjVZePU1bcPGtPsUI8KiuDmpiJq9FODA
TqEx9yH0MN+Zp7/MYCYgG/oyVdl0qP/ZA8e0tovccmqsBL8WPC2I+MGekSZWZd1XsQqmli+UNaUV
GMQqDsB85tQokDkhkkMDmot+WwVKAofUF17pP06SyCgkPG+aOjquYgKYaA+sh5Y9+rin93m+SRec
KaD0QNbO0qxJs/i/Y3wBnnIG6gihwl+5kPxkc3YOGfa4kNXcOWnQ8dEPvwXTYvj+aJOM/l+j3qcj
sNW75pRaDLA+2eiMWJxyXofGZzQPH/pbs5ZH/d8JRTlbnw9CV3Akoa7cA5bit1EokE/RsMLdbTFq
kpaQCOp2eIi+RLNc40A/B7DE0QX06xmrlpoiKlYXi3IEf1eEs5hIv8DNcwuempIYOL5SpnspcoJA
zl8WCnVwgLtQ2URLSeW+ufk0KEDh3qxgz1jH1dU8b0qXuJhCkhBXGRvyCD/1fvKcNWlZoL1ciTE+
IarXMw2sFLa1YqQ2VooEv3DIrpxWmBmF2auhtBaIphJ6suTQMi1QgKNeLcqbeRd+cxtlTZEHKVP4
PRxAKGQlbAtYQXbWAEkVkacBvDSOq9mkuyj+tMH8EIPO0Se8j6VEgfTxu/gxyaexnE4e4TsSWGXI
rwY4+J6lXgX86enOlQTSQBplnRS6Hirgf3A58VD+TpY2aRmjpEk0ks31fMRBs0JhyY6YzSesd+T7
NSRVEPNZ/8ULgFdEIGcrhnjBAlqZgsZi7D+MqGof9xlY8y01+bEaZRTlyH8ln7nZ7GA+mf4gOHEh
41oG5VWzZqkbu3aLVPJaqAibZtHewwCmx6Ii7uRkX/gAE7Ucmjk+TlF2ZpASay+iKX3SwGm5bi4/
cNYnZmTFE6dSajMMiu6Mrh3Ycpzn1q+JYEIB2Uw7VWbxyNryQQAi3B7/dFdty+yH9zuP6Qk926K7
ncz4eqrE95HfLZnvaHSIXJTTcOK0QZUkeF+NlqIfYp1i/Nmr00xoWVgpMgOhqJNNWrsalSkRxPNd
WN3gCVru4HDvzgrG8+IyM7VE+LzoM73aiGhSWNbz4uZI1/XO6R4zrmM5CpiZsAsB7JEt5HuE27OS
oQKpsFW130PuwIxAADxW3fI7/oUCrOZBaPOW4oI/LyTXGscmdgccEvpAGrrLgNVcmZ6Pvvz2nSaw
GRerN4ikfn2pSO+cSWsY4rIUprhuY4TYVsInXRvzL0Wvx0D8Y71zDGWVdN4pVKLHlEWfJ7UMSDX1
F4FyHi/0jeZK+kAEOwNIRuD+QGXqJDpZBJ90L4ENtEkCcpnck1IkhAXpZcTnf4FjqLR/91ZqMC+8
J2689Md+SMozL63cc4XulM6/LFzjPAPsfJVV8KgGmHaPXtVet0pA4jh3bGKcee986SlMCiRDNQ/x
cRylBt6q6riyMGYExmPHHi0OQGdPhErzxOJ0KV+LaG6Po5tSgXc3EBrwl1G5k/ZGdDWqPkCnmXIf
nSmniELRY4V4cnthyKp6B/nhPHThblvnVVaBDhWDBraVVyenHn/81EE6JoodnsfLQBAEdidr1Ue0
9+um+OP2A/8GZTrDoVoPF0NEQPd5RA0F+Dz7tRwrazRkWvp/cKzTnjHYiiC51Ubb12kUz50jKyCY
i0ZSI3zzGhH3GWZa1OOTOqPgmw/VIYwQEUMMbDPfRl/RPqsgBBET5PIyUY5xj0s7olbTcQMlkTDP
8GVJwt+Z8mW2Jd5o7+zx/pqhKSxb+Ivy3gKfAqmlhH5ze/Nn5TxYewzxNRK2UhJOpkjSv84o4kgU
XjzBrgn3swkA04gLKPGNflDexixY8S1+fcWflCYWdQQeogvV0Jk688priA7DFIpXi0jUXk305tma
bI6iTZnbFV7nm0pKycfkaCbT/YYN348roS/humwkFjOP7Fg4i6dBeRGXtxK5OG24d17G6KZwjifc
OLyJlBsQx4gB8+yMcDiQrNFM2TpcXyx+m9dZJHQmRSpGCUPXkcvN8k4Us7h2czRuvbkdVVOXBHJI
mTlTNxTf+tlhfpgKTuYt6T0n3HcXOFEEwXwBY3eB6zbpVY2vCfpenK7QcM0icfgzQ73o6Ed4ppPm
ko1oTu0/lZ5JbbePKjBNOPKSyftyX76KcP1rMZbFVXd4b83xZTBsD+9wLiIvQeZ/fAUzBl8rrH0Z
uuUF4uhAWB63fhUGxnqLcubhmH9QzwihILpMbePBfWqYKfZESy9ni5boSsAMcCuTRIlDtTXubg6T
sKtW7X0t03EWCgr8nDo7rCU9GQgy8vsvOIJcp97soFPFZcv3RMCMsomI0b2ftVoMmqWv9z2Vn6ST
0XyoUx7TVQRleTb85xhQ3djHrjy+HXGK3SoyqqSblUZ2n6S3pplP8v8MabyWHJfcFLXESeueYlVM
yQpTkTqx2QIMpFL81xkrNiGqlDKg+XOcyxNYBthw/mOuHjK4NgiCDPIknqV0KgJBwurJuLa00QMi
SdM3Xrc263EwO9pntd6W1H9Z4e/HZiGM7MjL0rWxurLCuok6bhzZsiB3PD1JThk0m463IvGFxwGA
tbsHVq3FmCMlZwvLVtizQDBPVLfuwLwBTR2Lc/IAEWIRqITgKhbl2Y2z3aI39Z7sktLgTp5tt8Cx
CS0lgwsBMYVe+89bA8f1EO/DoOcBYDNpab1foQ0mhJk+ZB2Oky8z+dQEH0xq3W8BvNKuG8ocG4YF
MKJToDuPDlPfWEcm4JnAtFP2JST6kxtX8UXT19Nn4ygWVHtXGiWfiStNlamTua8I9M/vf3tFTiD6
edlHNSWXgnC4ZJpHiOI6nc7L7fgDSlVYeBAlsX5g27OmyR1D8gEl0epsgwQBYsTfUgF+9Ju3ImiL
szG0pNKgFAvWxQAAYJ9Fn0MpVHl+fzBskiJdLHZI9tluuPTkQw1KDMjZO6OQs0TwypyzBAj4uUXi
QhOc/gQKKJAyQYPGCxfIK1UyQlH+iTIIpTBNcgXWaqIh6HI4kEwLbhfDzat+qE3aR8d2YDqMzp1G
v/hxUaYtMEbH5ymamHoYFTslTBLwtB/cm+Fx+BUngtGTz1FchK/NdWKcpeTDamwoQ0c74FggEu+N
8q7yY8D8bIRejZc4+RFTJlsIA0fTAd1mk1Di+JN9prPUhxXel5uHoNt4v/5uyWqgLjupJPPnvbm6
B12Yn6kFNpEa1a9n/NHcljI09PER8ESXH/3GCU/tIGhpjbLMWy9Agx87DfFw2lW5o/a6M/DfK9Qo
TYjUmctH0MF1lTrlqYT0uBKrdWk7p1X4O8ZvOMjiyI+Sqkfnv7EYli2W6/PgvV5R1zdbPwPcshrg
lUsmLeLMGu4F+6YmZkAmG+FCs7eN8QzEoIRWx4axMUGrkQ//N0TxeCXGVN4y5r6K6gXbBs2p46Ky
DEnpR02Lz5lCYZBViX5h8Ssi3I7J1th8UEasuCpPHrBt/x8JHqxWzeJT2ma7T6BbIhEM21Ji7c+V
qDJIAvcqG+3N2BT/mueH3flcte90fez66GMoYdpkirSHiL11Wt+6ZON7yqIUg1tPDF93cPevBHrX
kGJdH8eYqZQLp4yO8tC5OCBCaUUOjqKuiyVDlB2R4FPbYnvfnuEzxFAoXcVRxJke/LjssZ/YeFcu
nqluCrzEYN+0W0JiMFcELIu7lGUym87u7fd4JThssELsYAdWqCRNyro9swpaoJgG7o2gR55C0FNw
7PZuQrBENkx0U2+h1v1CHXeOMX23aMbUpOtKmkCm5gAyhcQZs5ZoQWJgwqGraYpHFJDjiRd7+51y
DR7Dw/7mqfMH/PszD3w07O8Lml0UU9BHR7o/kPEIWSKAyySs8Jj/Jp+23zc/pBrNKTJU6wdcMonr
PXreUmvkWCoVS0p1wWUUliBLojoGCDmj2miRW4dh447e2XOaiiHrrjXC7HQsaB1cnummG+cO0q+r
YitlHlMHukvKpB+qKqyXFQVwhKqdGNhrS/1gKv9yaJQD23UFWR4sRYdVfTmLPNFwI8gwkAVX3EJO
E7+4HovydEjEmKi92jWVjJyB4RwW7TfzaM8CmJ1/aPAFQkrHNl1t+2eoFRKeCgYxG+K///PtLn43
QhAHXPDc1PNwJ1evs6vBpcw1Td3sedm9pnDi+Xq9E6t/csDIIP70pcdVfT9nY6Q+Q970wIc4+327
TT4aWTvbboOmokkTZy5OxG0ygqOHtN4Y10vyyl25obvOw4eI6PEIIUMjyworbfRdjmIVzaIdblDW
YfZn3vUMjvKOsAijS2MD7oXSlPfRcwnEOdkHJgI7nXRy9obZmTvVsFrLcFPXt+JyezfoyXx5YBZA
bEG1mi/7mczv5eOs8jqON7dZGRIhs2x+3x68tzxsNIfnsd5vcevb0FBJpX4Mfun5R3zJNSVzH2mm
V65B5h2fzD2clhZSmLCow/45XUnvTilXXKmKL17/bYlARS+8lqPz5xvOVS+j7S1h9qYHft/NYgan
4lJ/ONnX6lfuQWCenucYnpGTvJhCsocndttmewgZuJlUJ8voOdckoFI7ZfMD3FlvpofZEUf1ROY5
YCAzG3AVLdvvcVRTj1uYGYMWtKnokAchLkiS7U4lH8dro6naSsvSChOPBEYGdlDiBeVn8nYbvvOS
xS4JQP/xq4HXXjfYkbxQdda+bhK5E2qh5N6Jz6eOhEcyAORWi3D86B4mqeM+/1Bt6CgiFp6d+2uI
zSI1zD4SBdywPO8g48R1PjZGoKggoA73YyOjjt377I6qT47NhEZ/hk+Am7wpDdRvTBrCiNj2Ibnk
AxIL+j2QmHEYUpHaL6xBNevxxUevtikebh946yP+Q4BEmyUTDh9aAo1fgQMpSx+fn+BuABx/VVYf
W6Jk21XxYe5dWy5/ELvq92jeVrmmSvGuWiJ026Q3v6D+cc0+7EWJEncuQpTpoz0n37MFW5aEfNKH
7JpaUnQOmb5EfwM1U4Uv5zJfwTPCGISRomp1csz7gz6RIsvatQhyIsfIuWyoJvYLAHr31G7BpCoq
ghCIgI6J7Z0YE5a6oFJpVlFze15fdCaFbwnWEBBHDEdNjoWR4C1FYv9y0Bxj/oG6yXSo3eNY7uf0
QQ4m9JVoERD7Vzs1Efa87RlLyAf4eqUf2IUCLpyQnEkC1pnvudvRd/OzV9Uhn5vu8iRfNQTRFWG0
F00jIYzyS37Hgnxus1G7YbJ3h0M0GLTeaachO20aLhiypge5j/c9+TE+UPMlALPdMRXsHR0xtrJy
Z3p/OdpBQF852yvksLbzCAiQ7QVwDFMU3PyTSh2X8XYBGGZAuHFIMaO+u3uHRE9a4VJ0Ziaitt0I
li6gORpBgsVxQYjh54GMrQqEChQrJEnmgE6BpNbQaPv00nO0AQazg7NMYpaaTB4n5YeCMQiozYIc
3AHFN6zA5GfFzyqq7xO2/z5IaBaiL7a34mgpEmbrMoLKxQplporjY9qf6mHNLkbPvfYoUC6uT4aq
22ibRuaTzv/Z1PxqDW+Z/JrOHCLxBuRB3npwAZftHSmoFPAnk/y6KAbWRTBYTiVsU7irzvBbbJms
WyT21xPoe4tgp6WRPmMgvhz1lGedJI8cripDUsJA8tp27H1P5UBWDrSc93KysJWvH19y9rxWrtii
EBV9NRaylMBEF4aQOWTJXqxWPk0F3nEkpRnJuvWVsDWaSia80XTrNiwn1sWhaukf4fhk+i6wFRgl
VUspCPMABXzhW8RgfZIZrwvzVlvMLc9UTttV3SN3miSevGemvlGaUevg6cjggA66T3Gd6ISil5X7
xSJe1u/Y7oDIlhWESR+tDrQbJ8FBp/fTCKyd+O0XsR/v7mjwR+LonumeEGYGgzzYw59gPPnSdXZa
BGMG5ZSoS4cieP099WtflQJcYK1reKHphDGSl0oZq+zbWfSJ4qTS38ImMF4JmZjQm8ILoB4uiPGZ
6CTRRxEBrsnjwQGufehsLB8e6JvLQo+Q8rvpjI/bRs/R5qoLq/PABEVY08mmQjbnTf+aV3gwIYe+
8wobtaGkUeQWSPf8C/eOqqLnQelvWncfR1fom1BHYJdGJlpnK0Ddwj+NIfLE+nXyrG3q2j/R7Nfs
SVD0ASOWy0EdyKt4CMxczwVcD9+XImPveOAhLh3oVqm997wfhdU9HcZrOF34BWCno8D0Ot/nPS9u
KyA4Zqi9iaYt7TGT5EN25SaeeWQrxYc0FFBs7S4DhVZDRt2vqgQenNWSyu9GixEDKUVlYalp4MtR
28SuMa4YZdP0KsEVbEQf1X1aVv3/SjHLAGoe0oshp8rFFlLnI5bQjfnjAtbUP1aozUdDgwZlmV8R
uMMzk6XEe2XP8VKMNef2Lbjo4aXkVL3e2CiPvpBs6o3Yr8tM2Usqp82ePHG0YvtSoeY411by3DlN
mrub4d+UHGDrJ66sZDJ7N7iDkJbwjwpViV+DINHAZTK7WUpMf9jeRYUzTfb4nQPjWO9N3vHsvQqh
7nyLzU7NhRcuemPUHrPDkHZDE02iLRENWGNdHLTj9fuxv2sO3OWsntxxvnBgbFedySkEIm0Nuxey
X55NWJf7OAwV/jdhj10ZcYhlaWaKuHvWHybs5rZaFA4z8Yl1+un1HH5poiXdfWeLbPF+vfUeqKjf
6+prdJoaqmI3hg9yGk9gNkqC+X2ar7+yumv8h/19fCXrXbRtuce8nPZGJp08QAFMGuJndMhmadE6
W0LtsM/vPkM+Mm/bqT8p1AEmFBrjGZ7RQmMLWlCRPLpB9gMWejXRrg5VV+DL9Jmb/PHhzrW/mEsB
dt0OMHp3utj2OIcWHcfVQ7nfWbegR4rkP4p8WM9RsLWRfvEGEsGGNlKjM1+evKM26eBZUlar85nK
Yp6murMpWa9Xodo+478idtl7xYsVWyP1hPB8SMznHi0W4fB1rZoSe/W7ytisKxGx8mtGujKQAHR2
p1B2zRcOZjJawqaDzd5FrDdXyaXO4eOQ+uUbfQ8x+VgERUrlKBaOoz/TTa4luVk+SYBEijd4pi33
sn2F3FZnx4Gr4+E4nZxdRRwSVF5hH4Rmk0fjO/2JmJuFJwivdWUqWgukBzFu65edqV79PU4H1PIx
a++Q5MvMSWvpPXUDCJDY54VvwjlDHpMMlEMOwj943fmj4JxpXh8fj2BNiRzjG08pvYkNUKhCVzpt
z0a6+azXQL4TVbl6JFwFJTyy/L8wlB3al9Y01ETNY4DVjgvb8TgA1tHvD+ShLaGs7ujJmiqyxxnu
Sv+E/O05a8b0XtCJq1ZA2Nva9Xfe89QUdiaYfpWnoqQTkRF+dGw5sfo27ifKh4F3Etz715gDIikA
me9W9LkHA/sK2Zstw9mgqcIJZ3hO9giiwtv1epq3zxjLpLLfRv6biwrrGZJ7K/oPGwuEem+O6+qT
PycdpVx0KdsHSwVVKrjjIwt0oSxPqqcFLuZBO9LP319B84t/0x9wXzDVyMjLLXEeV6L1neJhVbI8
aFulTq/F1uuiOhB9A4kFNbWgX12Ei44lEXFvi4o7wttihkUJJGl/NIQ55tzcOoOkvDbYqXwSXhMY
abmNka8mU5Zu5i1iPjN+IxynDaq1j/bSVKXLoyr5KL3Yioe9QX4nVME4YJBHHMh8zHroueXh1f4w
6RDggjT6Yd0ePcayo3qAcqC26+YQ81yDM8wQv1V079zi19gf6KJNW67SECfCetsRmy08ABA3C1+M
yROUyKUhwruhAYaWUVNNqva079umAQy9BwJRCF4gZEMH3vLBE7pKV/8XbUSW8PCOxND7+e+vlGjc
heVZWzURN+MgUPqZC2TbnDbmyjNhtVcnnvAra+Takc3VC0GoXM77kIhZCwewLY10lfpARWnxV2VQ
iiKBw1f3EeFOVPo50v/+LxJQE88JXEssfyoGIb9vVXzW4wSHMF1BihkWuQJ1B1HbA15EwNBNEVJ+
8zZqVKgPIrazL/Sopgj/+BrCBpTr4eu3J4U0WKc26e9wQTbaY3j6tpAtHCU02jvRiij5LY3+T6gd
NUAxQ7zGDC8akHPzdrtA01KXVJtNg2DjGrEIL34uSoexdmwfRFaLo5yZ5Gm8jIoM/sPjE8G/Z2K8
IDoHKU9c+TT2Tiyx+1gfT91+9YOylAXD/WXRfhWMDyJUqjL+iG34ftnCT5ZJNHkwR+WDBm8kQmJ7
DNhvN9D78g6+LAIsM1OHRwqyLbxAGVih8SqnVlm08xN9sKjmB8A87XvCciHxCUqqskTELRYmA1Tz
Jt5sSb2o4uyrbfaaL5h8JfhVZjZSdKzR6WFY/HWjCo+hfXgnZq6RdZJoX9J3OZFrKP1Yc5wNsGuK
WKgGYvJRrk4sGfNyMP5XEbA8KnzHlst6UkzeUnFSqkmUIcNWe0AsyECD6uhJYn1D2lrS8tvsoc40
ggVTz2Gn53R+ExYUgi5Sf4s7bypl9MYuqz7sXpStg0hkx+EySlbkkaa6GWCJK+hFNS/opLjDYkFr
vaVcZ93gEe6BzvGJJQaziDRWbWP0Wygu8gtkNnnFhx06jZv8aSj/vOn1SDf2IkDRTJ8yHXGG5pdC
/JIH5CWbVv/k8oSTSHyHGzNEHVzPERkomRGCNhbA6Qyf7mk3oRAArFRjiVi1fqPLUJcT7bQyQFM7
G4r4xCZBDsD5VsDecCfN3uH2bjOnIfUNOe0gw/mE8MgCV8kO9Yaz+7aa8en+ixMD5nTiM3E2Lmsf
7fFoDCgXZyyupogYZBHzckLPdJ0dmarSEiETbeN3IkU6oSxqBeA6iBd1Hcw08Wkn/X5UTG3EqApn
UiVBdn8ATR0BbX/imE/oh4aJcB6vHi3Bq1v6DusnCnvAqlES6kYn1Wog/TgBOo5J1Wfsis4wXg5B
+U908+p5DKS/lvCK/v3ZMADlEmLgq1akysTdp/1IaNsaDBREND3nal1YDmkzMNQFEE5aHI/YjDWf
hHyBjDvxHJ96pcZNzaqn2Jf+IgfBSQ+FUH6a+K0c8ccj1ZktqotWzU3D4SnzOmdjBXJBfkROZ/Jx
Hp/tUKOIFMEVF7Zn4xri/8OIFeW30P066g2UfHks9/F9v9lde6pKNeFhoXirKDLtgSG7XqMVgYue
JOXKqcvnPDd/RZyLKvfbchoCqdr38/xMjTT0AJYp80CIBMcuLgEVAd/GkqKEKi30BGSrgPHqaJZ3
Z4G8gpwCl2o1r1RdtGY+5xzGwkN9LbQrjh4A4L0tWSCIbujUXwLNNTb4L/p9yLZQfiiLxmh/kRhk
2sr/2oIiHnSjjq4NkAxzehBUYHY4bVbbp/zsK0wynUBpyyIat+HdkefdPimRnjyrQOAK0W0s4J0P
9amWbGNsukv3zYUb3+OIReiDRMEOJ2xKmmEgtqdGVPNuXhOxB9OLFleKavUT5TLN569M4Zwt4m4w
M1fcO93NzoTmMqKUlj8/KMmtp6nO+qaWoPDHb48Js6XRWhhcllvgSrRKrSZJo5vZVE+/gteSKmZb
FtjhUGkZ0jKlIRqfWYJ3KiLEMNozSjwi92JmJRfBEcMSfjOtDSPNsOpsQk7K3FYX1U6It8Vnm5eU
8ELHeTfaGeQHgO94MxfEifQWdwF63d/WKb7zSRWvgDzfCceBhWJuXXe2vfbXc7OBhLxdTnVp678/
bIhLpXgrxwGmtbv1O9q0rl16CTmwjyvMq1XFoeAt81cfWE15h8iWSM8eYRIV/HGc/NWLdhO9y8ac
+ktl8F9cG0Sz4hNEI99n7Uu5T6Zf1Esou6ySdMvUL3r7pWtvy9+g5DgaVMC0eVSAJodlnwOsQ3SR
dTu7sGUivDSYgh1Y4EfrczfqY27KbG2SgcwngyrEK31MHUrCoYkZ3P0nccprBcLubpEZTV3ztceb
arfD+j/v0qoFj+Uvnof4GNXzITD8/4mDofgGzbPn59nSeBJtESmKN8HodguKpQQCVxWneNWws4i3
s/KQ/QbYEudyEj7EkPuev322yiQVw5tRPIvZ6dBkO9ZsmfqRx58dZXsxFWKEBVETfUj2t3dS4Uhw
ZcooXgA1F8gwVfviarIlQewUuRNuFl0BKOItBClJLz2lqFJ+ey0XBFMh9v8n3VpqNvh3TsMaJOUd
oNQ9wbxc/JApSjxuRhMFDx2QniHRgmVGw8EtMWwfpXw19Cwnh7tQlO9zTr5Y2Hg6yYchXG8HmvoF
xYm4JtfSglTZ149ZFjZIfYjcl4NJc6LQdOhGeDKkI10NMU2MIU7D0SKMsiA/viupqWzF2yMoDShB
tkIJq5fupXyl/iEcwDpydPKfjFg3361q6ionnj+kx1m9UEoy1DQXI9dVoeAQFE0yQJpdnsy2MWHA
tkcLmYnQtc20sKPn3l7ykxpH+z8DxaIP+Q4xWZWZbu9M2SQZ3tm5f87+OGh1IEfhUHtfgjPdSqFC
Io5MsnrvcOFEjaMJV8B5FfUxeHC28w0MLEXZSVuJEIH1wwUJqMOiiaXTjcntN4UduFtXwq6Xd7GP
QmOE013W8fOOJoubP9fNYBSDlvCO79WaQmzNphUPQIJp4wcPyMrAKyokaIK9k+T2MzuOQfkCSwb2
bfjq/HBodq/aETAn94P3MNVWYeUoQbFi0d7ncw5b8evUIZlqMNOE/yiF0EjUNh5QoVRimRaWk1I/
4EsPDL/UTYOJZefELmPKFOcaPpa7VDSB6qYqavO8LCQytXppwfD8Sd2l+PiV7Nxj2+0pzD1GhsaV
iwG2KQvZXvPnTIR7c0rEGvHKjjG+ksiV+6GLJ03Z4/61QtPY+kQTpHFEhoWhVD3j36aRVqw7IWJ8
tFYN4q/SJSmZagjHytdZbQCnsX1a7FKQBSbFeNK0WTE9oS/z68L0ooJtnbv97ICKoxn40p+niQ9K
ssk4cb0iQcgfcEV0aNkXmMoUdxmHAIkG0JcQOd0sgVkph8Va28C+waeC2q06yMZtwdrwdNLhEWeL
i/U9OMFko1+Gjfk4UtYj8Uj4Z070Mz0M04kS8ibfj3lxmeSfLhAdl5rfiGIiCopFVM+GddtfA2Ub
zWBGg3cUkkQ0lAAwjSoG3auak9xf8JkpBUWnBkxXL7sSEcsqSFuYwvjJJTJhxrdqmd018RRPH9dL
TQYq5BAoAYNwF9KL3bmcB72FORGFhZj405lrpw6ch6J4KXFw+ULtr10SskMr5ou9Jnxf4u78Mq2l
kUd1aiNHr2ksn5dJ7fzztaNqkWjRq9go3Z+aw/UIORUUwF9WAVacf3lXlQp6UAWYnteqnxbU8qIr
4Zv/KkVcIxmlSBUbdvbfq9ocY5PYf6tE6+Zc3EG4IOaAlLFhit7+JZTFI9LybwDGs4Wal2X7HcdY
l07mWf9j9pF71KAEiNIKGS2M9VdNj1AsbVR2v2yJLEP3eDSgJI4QSGgL1PO8BN/Ov0/S1Shqf+4D
Xd09nd7GIh+kN6nyo+wuKczQi7gviNZyG8jcXhWoBGnMXsLWDetHteeoHeEuH7rMloXjpAJmHnxG
MMJibMWP9dagBLwPE3ZidSBWBfRDGBmMHDVQNi92xPtMazd/RvZu0ZnTTQxpb1azeCmqv+L49sCe
joBahv1ooLIbe3tIyCxGX4Y1jrJEBu004dETk31kIwUVgvFE22xVy0zpMbwVjIU+AgsJ+5JJTHPu
gvxglYI7wFJOXPZyvIR9KUXpTYG7tr+LM5B+OamYELSgqtx0pGGqvCuLZ/nN7kudRTLQrnIDUVcc
5LOQZ+d4bGN8K6sXEv7kEX3poEHoA0N2LybM4XJ1PHX4sWwupBeVrOfcbpU70D5BizQBgPeJqyiW
z6QFsGBNhf8A59oVXmbIK691u/J+ZvKCeukPqzAqv6IrsrBwVNUexINGrs1LffUiMi0eqpzMS3At
HozIbyvfnn8aSzbyrE2U2DjzUGoi90DcOtn4us1aGyl0OH7FCa6FQ0GVoIh7QEWz8xKRnDXISRk4
DkLTkAh8B3vdR249jvdFUaas4LZNYFcU6QJqQOyGLBlHl1epdaoI1BzXt9SLXzGh5L+OR/xyToOe
SatgIlIpaiO5R/SdqAbdrGx5JsfWqIa0lz7GmXVmw/nQdXmGUQaBwHeMLE5WxpMx7kmU3Z4+xb9u
mEpLMFg3sxnTKXVdNOyb8gYENKn0YEnfCeDpGdvKp3wKrCjX7e/lpyI4PZB+ivJxHn8r85uL5/mZ
m/2xHM2LtwujBp+gGAdCRnre7z5lfq3W8rW4cweLhiF8Qay9VS018VKF2Fe4Lw6GZenkhnnvk20a
wCJwDDiLk4x9w5RiyxVcspNEruRRnwm19Dm4hJPJtjdEJTv6k7w3DIZXA6NmTKi1+P9cobhMXWYa
cLEPnI1+2q6MxYJZJr19d9GhFn511khknboQtTkSTkTstL3TNpDCM1IVz+B0eMkHt1MzzUW5CALn
rn1Qg3F3a5yqPrRtBSuP8zVTAwKGvTid2Kq5ifXSpWDRD7ibJhkHZLIVBit60U/yYDL2wsoQEWXp
+VdioNMUoG/o6Z5xzx5myfdfN3wqWWeFy88oca/cAiNVd+b6hR3jiNYRCB9wUlkKKFMW4024fWXO
vfE2WnF99dNbbm9HfKugxAMKB1ZpVukcjn+F1yRW8NCrIedDCHfqwab0/9gmmvcaycxaLW03uqQm
krj+AsyeOT7T+abYV5+fKOv6e//zdyHiM4uLBJJSXJao1zUHGwvqhaqjjHqc0UUFKqbVPIDsOD8f
Vgowv8sm9Don5uwqo41xuibE+6nowzioi7yx5OdAcP4pi4TNY9Hh2ep/MESy6i2iyV9VhE8aNPdz
P08kTAfS668nqfhKoyfdLSEwsiu74T43dfmiDHeiYkcq7v3X5sFmpSKpY0MFXKQnGNSkbbIc6nCH
LFbj6ELkwINLbDoaaCoB7JcXSgbMZXM1NhAIMr3XYpTQU7fWClHEEmDdNaCclfYbLw1yN72T5sRT
6whOwyhx4pQOKNRJNIsh7lJW2JW/oZYE9JRJF8TYE9oO8mP5W24XcmdCr8PIwfMJ/cMCdHXh1QxS
0d4GSGCgDpri+cwEIg2+O0AL+JgbDhiIB9k+F3/59jbGqkEUZZbrnGT5BBcfYwhgf23eJPeBcShw
rFEBwxb8hJ6BQKqM0N2eQMyyyEpY5cVEeIQnKTYi7bJaC/D7RkDcVMl7U+1okwea+FBubp3kwoRy
9+Ojbf04HycKeic2zlEJeKLsyMv7AWI74c5o54h+qOrWbFRTa8hm0tcWhl9Q2dbalZDG7ytAkZWC
+anMBx+oKD5tEctb8SVlePtu6FwMrDuskU6kQz/HBTgLat+Mjp9Mnrovk8UKHQwpjUfMAqQItHel
/uJ+oDsKh/Xr36h4xovipY9+kDFNMQmfXE1G3WNuTjXDFUYD0zD0StBKdwwy+QzluvPqg1RKgKVM
QKaFALJsNlsv5ccLlNeivXvHZlOqdTyuqTlBKBrVMwSb5tk7vCJ2CazDZ7T3nBebEkSqy1bnw2Y/
qcWFg0ZV3dvESCAlZtN5edlsVTg3uao9T5R9ScBeY+iFOctSt0Ycg2i2fb1nEnTUO/1Nqv8dPNH9
Wy9Xh0vfcVM/yVOnJnmklCKAZ9VoV/NYHfegVY4Bj8p4tSgJBeIcLchOUMR8XectYu7mACXwXDFz
wGrHZkjZMZQT6bsrZhxcZ7gAznrLX0XzchCwGFxLi8uNP6OvXVmjiBEdxg+kAu+JPllx0nxJr4tb
Rp1LpnO5W7NeLsADd9aOnQs8URW5OZlUvMVRIOVkgweMuWIblHuUAX+tic2hHrBsSQ617fMBQeM5
eurMF5wCG3cQYD9xJeyz5ddYvPtoBAyjxbb7pUted79cCdWBRrpPxMphjBUldx+MYEbMMxBgHwoi
1iSQ5KsUaKsYIT25KRW3Xr3Xm8DR7EOtep9d2531xnoLuP/IkwSZ7gF+P7x8srV9uNZkHtf18LA0
qm+sBhDrVH2g5Dbhlhng+cCD7q0uaUQqn9a+yB1/Z+MmTsz5kmUxV6D/bRXMQ9RR6dfejMMzou46
DJvaJWygRzJWXfi/x2skz7/c0rMgmmjvqEqJIfhqEHaKjxnHdftZ25gX+KdmBYiypDuvgI15Xv1e
mhsItiEEyXySObXjDzt/9RfV1orHjbXA/Vc44TK+sUppVo/gsBbAy+/nG0TdxJFloUIwCpBcbHLX
tHokSYnjjm5XShLqfFn5m4+Xer65JBkYP2zzVqYJvjhPFzJglUnSIJJ6K6kSL5xyKUweY5Xb5zrd
Ck0T+5vVrNUuzu2HWhEVfH3EzlE2MXmBObiA1QTinPYrXbiEgp1WH36oSWHYLRvbO06eE+vaAR1J
884Ud2GCdKV1WzmdLsBPo5zR9hX/K3RAtLdnvDhv9XrRvW0YCDmLwcU0X78ipOQz/N5w4j5V5Eyb
q/QgN2rsQ5q4gEZ5WEyCzSXTQJA0WebIEoAToGxMTlL/khbQ+IeRfOSiy8vlG58MqnyHjXLu2ApC
apN6DVjdCXinhgH28Z3wscKsremt1pkRpkxoXHSHHe2AntiDG/kFs89Sq2gTxdO2PB2pJbwJiDJz
QuliDCIFuz8TehWlpb2471SA+2Z6lMbtDFYOBj72w4MXGWfxVg5YQqLV4H+nMYCc9/ePQVJhWx8v
fiHgS1WXG+RrNt7AytApLthhXRapO9uT/p/eEIzm16kU8x1qsLQfv70xBc3GnX0ow+4Wd+euzE5/
iVQXnPsnq7R63wUPV5W6dh6EiiVkf8ODY5kWmclwZaY+kU4FXka0zyJJnOFg+DVRu7MFlXFT60cb
ALSNJP5J80Dlc7edCJk0UsQQ077uBGFAC6TAXnqjCg7/tnbHPSwK+yoN2NV3O+95kTjX1hwD7WX0
dFnpxW90UccrSzkr4UyvS7i6kpa/175001YAvrxe1UEu5LyEG4pEkTfl6b6Wk2klmsyYy5UBQ1cm
G0btgzNG2crc2Zr1qUaPKkC5Bg+DkqMPTS5exIP5eEtHykz2Uygu0T/1OJEUDh63lPYwuEor40Bj
QFPxjZTrkeaLAW3/Ablblat1kMayQkME2q4ElXi5G1ljBLpForW5uxHdsMQx1UR20++cLr5K921K
9lQQDgJLvAj0SnS/zkyK+YNRMcQvbnnEaVciuqnLMgOomMPMqPrcuLEhyqjX7skS+jW+o3YsFVIL
Regx9jhzon1LR+7kQg8hx0X3qEirlUXrpiIBd3Wp7IDZErnxiCuPMjD6fdThCNg1Df7YR2sy7s1H
JdVpc9y5nfn6bIuNi5xQevcSh6/GTxdhtKvlSCjp7UIv/WVYe4Yz3kXbyWXBTjja33PjkGyE71M7
+h/E1Hkl4adBst6fbfEIIJkmYyvH/8oH42jC1sVuLrAn9OdM4GYfiMQZOCkuYN4LUazcCxD3e8eX
1asZxPNC1+qL2EQzSgmH16RNTUgy6adiamQY7TVj8egjE1mxQiMn4O725KBS1bSJh+fTHh+fIAJd
bvWRFPmGSphXsiCOWJ0EW6V9cB/TreXEkgam2ihDia/9OcDcl4Zdqz/QmRAqyZ1D0X/AK3HH9bCj
3ZSf8LbY3WTdZVwg88/3aCCkeRfqWC34MFo646b81BAGZgtvH3EheaUA90tDrOgohTKN1p9i4aYk
fP2w7yBG4U4UP1BSmT8ACPmYcUIVl/QEd/Enf5HVgXx7wgdochlAfqtRrABAVO+CnJE+fWpRaj4A
x0rKvywAW8nAMTJgkmLMsGesWklRxpvE4n7gBmseQxRetE9rCSiLIRrOFALo4bmgbkAqfPx/983q
sXP9wMfZzFZMjbm/2YdQMsMnzc9IIbPSqnAGcxlInGBVHWJovRE2EUsk0JcWJ0M1swiFc95Ec8o8
vNF9o5pq7LTIg+x7bVJwr4YdHi86MaareNM4beIc4w1EiiZI78OjXEEGYWoFSs6vQCaoH1NGQ8KO
Avo0hWGAvR3opTz1opKcAotjrb/SpQQVKouHWbMSH4C3VNvx/K24tfJcOyXI67rLdBKb4rc1V5NN
1NHxl6vdi9o8MFuiwODZp+fBvU1CPGEr9th8loDAwmn7wd61aGayP0YiIg7VrghBWif5B6TQEjeM
DeRQ6zh1gHQJPjzapd6JsbSiNI0Il4PzQdJ769ke8tGUlWEmMy1B/eUfVrtl0i0pfCaLNFEph9t8
ksKdC3fBT2fIO2i5zaIcpevHFhN/IJraJihJelFe1YdqyQD7kpCYkeNnWRtvdQjdp7rTGsM4Qhk8
iEGY80B0eMQhtYn+OLpToeqZtnE1MRfdsQG6OaVVUgCoqrEd8rsvtH7W84pmapKCDH5DK4SiAieF
OEnMv+M4iT8vsxriCpTgU4eq9TKazbEZtCzuVi0NuFrKA06kvuWMphY7doQygCpOHp7uz4wdlTp2
apm+XBIAivIr4iPWaZ6ETUFtFHF4C4U1QYBomblbX57gy0/c8kGPnUMCX7QEV7XVnCtPZyEPSU7p
tF34WzjNxP2Cv3TMzeB3kMKwc4uyasZl/IgiCwX024165rNHOp5PgIpvm7UsvSmTUw5Ka7Zuddr/
7ZtKrJ6l0nxj/VJ96GZxEg8pcMrVtkaj6OX1Cz9vEt73KWjC7Tkayfnfy4Yxd1clwi+3fnCzYV9b
/aiB9JQpg0OkoSWkwDOfWhMKG1dZOhEpJ88MUqR5Yy8FVUkZlTgQTaWdJmbNrHmbstdRw2Xf65X3
xIe5lRuWUjEtlZT6Rd2DrAhs+ZBytKHlsGTtMCUgloE6AQY7azQAdic62o45HZjvfrHeFqxKOYOi
+9y/4ZHIL97Zl31Z+0XcQYpxaB3ReAoBJy+iGjc6Xiu8ipMNVQbH+lrCCqQcyvQVRaN3c1cREZvj
6+mKkEyeq7mDKrrhbmcQ+wLArzBrP/97dRYne3vwhLW0AFOSoAivHOdvpUVp8l/K4+InfCZzWVLJ
+gGvSArbAgQAFxglZKGoADWZ3HxfqZ3fTh8W7VjiN7fgkxZsABPg7ViuJTuDpTvicJV0CulRu5SG
7kwCscDNO2Y+pnlOcP+sKfjRJBqEJy+fPY07htJY/6vXDzKUnC7KAGtAX5TTOY41MhQ6IBX9mWlh
5poQE4oXjayBBmpNrxVr8/tqlqT54X/ZRyMUptzW6GlvacnmD8Fbjn8aoB0ZR4dFI09ZXkK0bovA
MOTooP7F+3g+L9MLOqqjft+bABHNftLM6vvG1IUXARmPZl17Si1rRfSgIr/s1/yvApYDzqhNp8WS
0CtlWejBZ/OoZkIBoIzAsAWU3osEttT5B+4Hpv/eI5DgWH+An23qgiksx08wbEZ4g06PRL9bkw5Z
694SbXzP/2oqd9AwSF6W23e0JoRVUYLWZauqC+IWjvD+L1vxzM/sz9pwoiu1OH51DEGB8E/7oH9E
PUGE74NfzvPwSPqhMfiNBEpPCpGNXhxkH9LUIV/ewdg+rCBIuxKs6clgiHzUV4sHObX5wam3oain
xQJItVx7rNnqhILxYpm5V4T+3g3LfZ+7WNYlOY/C0kLEDkhDtIFfRFX2SxJI2mkS1ACqBpcBCsBy
vKVxbrStKohnkwnS8IgNMjNUKOZ3HES03yzNZoYxesTCzZb7dF1wHdAjdxS+KV0wdQaP5xchURqg
wKcZMn8822ikWAJEFklytuSA+pgUjXZpqyFBsXQHCTjM/Dx+CuiU6wXqE7yRuIkTzOm5+2sPoc1f
8Mnjrz1/hwPnS83r+9xoQSVx1oTEhUE8A1BW//rq01SWJOdS0H2JPiX5aALYjIafTRaSAIcv5EQG
o6ckXBpy4ZDAai6h9sffShV+GAwiOq91fLc3Fc1IThQwhORiPT7h6W2D6ebbJ//4RNLQVVdXvzHj
wc9nIUeds7qP5zJhOnGcaQ4k94A3bI3K1tCzIB4rzS4lNjoXadD+MvI3Hy214y0iV69+4Nf8dB3O
8iodYdrMByUI1SiD4iqQjeQy3bwQaD0cfYIuEULUklXLJJbvH9RX+Jyp+ivwizQBDC/Ul2zvtaNG
zqo0QvdnQ0Y8J9tjn2uB3eJ1QElMe8/CEJHz/NvIyB7w8gXpwvezObX54AZH7DPeskOr0FvJvCpK
XNWF4X2aQ4MzoudPuF575ms1jOHB2+HEhfmwXrT1M/Y5+qS1pBKkQwWQuyXUrc8di+qjdo2gXLU8
RQhHfYPj21VHqlQ7BsQ722+lcNVcz7GtznZzxKKyt8NX8o7wMMTtbptbYslT5xrLQZiBavOc8zbJ
pBefVLHIVq67hiZIPijcQvNnyP20jf5ugqZ8QSqLT9pyHLEaHa85SeqAjdXHyzqP7nC3n/6bsqPE
7HOEAHv4s+HQuCUUI++Rq2BJsqDFSBbDVmAkjnMAxUMNXAPiBXsXAFePrbX8Fa7xTw3nQJjF1AZO
aiDFjNy7jqJSbNkHHz1V2vXiZA40D8t/n1xRBXwJgNVCXmxVsJZCApqEiGhQ+UFyEEdDRLcuGVgv
L2PhXZMgtphSJInGTobUkB/ydGpHKjnBVePfVoVJNy2SFpveFKQjL6YEbMg/vbSlJ+kVwWPvIpi7
0f/1eEGR9c36/ZFrm3a97z7aLg+l1371ax21zmfROtpbtJGVLaufQIBuSZYxF/tfHigoWkT5hrm2
1HKS+AHAxwT/PnXItxC+ACzDc3thVloVJ2xdrFFb8uftuiEgQ5JdTHe1V0LK905Ku1bp3aS1jneV
xT+3/DnauQLqwl7fvK8VpHuGGMn7r6hhrEVgSjTWVcfo435ChX0ChcCdQOAZCAnY88oD0EZr4cOm
DohM54ozm+1GbhRVhd/vjecwRmDXH5caLazAdKITkP+C3uMkx4f5MgHW159AlnZlBsXDIU/dvS6D
QlWT6kjya+ejGfyVZPCX4YjtbGjME/9mplGSYNZQ8NdvGIOoXRAbA3P8A3G/y6GG2jyxMUUtDwHI
u5OvP5uwtEK4pmx4pTi8eByz1zBQ7kUoLzFIYJHMvJihkyy6Olhyc8yApPjC8M8yBOABxUwK9I/1
TbIIHT292zGdElW8SefJo0p06Yxw7oNuoQNgJ2HUEIGFGRBaYY5ZYIfG3jeZoEv/CvY0quvl8pFq
E0QJTVtHVnY/qaBA0HeITpx13ylurQg4bLMUYwbOGkyHqtUOgxd8OGu+XUMxBkwKcAOo6pJT8aR3
Abhvho+dHsatoYQGhZgMR41HZKvBLsvUZWl37g0AIeWf4NZpZEH0YlivmUZCLLHWFCXwblP8BElK
yJeQxPCkn/Q6sVzxearxEoap6tJHl1VUn+pSPfXXKIjNYEO9p/RBVEmyj8tmrHMquoz27RZ2scDo
JYiJgaLL8egR/Xo59PiI6O0OfCZNezzshBEiWyDPOq7BAP0d423rMbrNQCCKPUUKOmkMEA6vDqu9
96Wj8jyXAl09iOYJ2shVo0mYQPe58aAl2L7DwJgZj/tJe4FfPy2jyg9RH7mDLRbrE9B++UqiWZFM
peFXZZVGecxjNgtJb/zqFoiNj9X3EkAzm5bN7wwnKubx2iSpMXyR/jzA9APYcmsDVj9c3414RFmE
QtpaQWkfRibBCO3FhLKwmsbc1NxAduSsc/kpdCKU9zKV0V3Kki71JKKAmkt2vyg/FxUtzQLyQhfc
hMQnPaFNZgrEOm+bToAI70lIThpoztRl2+xoa1UITuncP0nkD1jU74bV7ph/0k5QxBbqI2R0HyjB
Hu6gIzj4vsPtjP0iuD4WrJ+4nhxtP61vSmyMti6WuTZ304cIMxoERbkgPtFH2RVmP5vOPfrbqurc
Y+CC5chu5jPf992BIDO7H/Pz2GCDyfrkUlt7t4zhhIOhW9FmZcPfwBPhQd3lHVczHbI1vqdViVvl
vb7pf76YrHpRwpJIiBKrDRuNobvF/0/BbwAj4BXy3X3hz5IWlawRK/LN2BfnHrHT9TVJ1Q7HU5h3
epWXFiK2kOiypOhvFVrjcUTdS832PXV8+aVWOLzMGlMWJG8X4q/boQgqqblRRKYYK5aSx5RgZMC3
rgeDXJtwLAkTKAqZvA1H/qzR3Qg00o+fmgd+hYJoIoeshmWGh0m/yl4ZRuifEE0/TiWmjaDVV0le
hmRS0FquK9YZI56f0HenPf188hkcw45VMy+CFFRQ13aNmxToY+bVwwQkWg6UVTBZNIW+acVojdgG
GpvQ+Tuv7AVUDUx2pW4ubJa+iOUfcORIhse7ONd3EhqkrajPqWdRGBl4i8Qpia7hhorRH0rkT8pm
PE/4WMuqVecInj3MCpqufQxwj91EoSkrV+oh5f+Hwceiwql+aF8IV823WUXQAz/WGTga5K4xAeDb
wihG6IBTP3R03/iNGpH1PqZfvbEow7Uz53KqAMFdm1zqG24lf0jjNd4edZmCh9RtViQriaThKSJa
P66/LGLt86yFAM81fPzRqckHkfA6o2WfrQFcEF0GvD+kGySGJbVMlk+fIg/h1AmyqSMbwHTBwfAw
t+aaLQkzxci+2XX4RL9xzpkXCGvJBQpMPVDOkXyDF0W0YyAU5riAcDHjuqQRNQN551CiMteyb8m+
j+Aa5HqUKlCmFLLzrRtRn9G8L5gt3fMi1amlpOZfuFPz/ISC/MrV6e2QctqORPLtqSOAOPYbM7Ee
9SM1C9c1NDY58Onhpsi6414tsvgVNvorqtCDEXs1pa/vuObYeLuLxKJL38GctvjTsINVUfskTojY
Of/UK3Lrz8gOS4AMWFO3mBPTCxpyHa1w7sJ9nmVdLMuxIEeGvdhnd4dvwj0aGGGTwKb06747PFzx
ceQtVTWLj8umuuVl+Y2wPWDZfMcMH/tp1veBtUzjiH/Ck0DoM/FRgmCaNQx+VHo3L0dkxr2WIhn9
pZ8h4TfWJ35VKu3abUoqN9OJB3I1wB1XsvcaT7hTXiKTvQVT5IaDZfbCq40c8CoqKqAlFcCTgnZC
QThSRGyI6HrkXz3ayxYOezp+mx0yuUhXiff3YLAXmHvDlz2KwPSwpi2ogAlxtsetiXlL/Lqzt960
f/sO3WwVBH15fvkZAmShg+700wWaHzzXR6xbopQrEi6W4LHUUAoUk0w6mAzo3fxCT5v5f6WJ9LsH
UL3IR6S4FgMbCQeU09Bnc8tNJPCN048Bo0QGYxABGwOkK7eD065GtJwGW7trQP5biRG1HV9+itx2
BD0SIP+HeWmNME1qjk18wkEMRiC8lAH1da+DaTJb8sjXLoX/8g3iJkpuYBJJAMSTjS3FBF1UjTFE
6sh4Xq+iPs3W46HvGYzxkNsDLvHmdYvahadOf60Iw8cy6s3B5dKCb7FWoAPY3/u2rgDfJrjdEafx
/vYUfUuaLs68UM8atkniZ3voBJqjXFIoBJ+cefMDEIELafxJvw6okhttwVaBf6t1oLIU+DPJ3jnf
Z+x6MzkaAx+N4Me0176zcoi85wN1KFAdXlHsbc7FI76Xn3oCRWkEm33ZUXnRGtCe1dVdb3/0XpmW
2ZQUoGdLuH0GmdMYHjOtjyKbYbpf2mpTRjyZqSuVfBJMR47CeBjSli9l7R/qkJwl+5VhKuKuOP3P
G+G7GrrpkxAw+dcSx8MiojDtLR45mqIL8x1jOur8hwdwQptrqSGrkbr1i6Sbqqb/mS42QcqnZ+eZ
3IbdDG5en5qad4vijd48S9jtBxN6vTG/DLSx+HcV0KsHlkJEHtR2B6Q0Mec1SPg1Lp+zXBXwJSTi
4ZouH38lGNYXshdIJ3jo5fhhkYu3RFygarvjjH6UdN3xgdSRUa6mAT8V244L4kwYzQ05xDotOJgy
bp+KmFKPYWadallUPqcXY5inz21ZhEuyvMuVDCq5Rsm7VkLJtmhhCxF3OMOhO4VhVGuqkMZkCBuu
tYQDK1V8xmLMcUNpAcrePlOhb7uJn+GhL872CuJ3WqpZXKLDyTROd/hqbIP1ib5Nx3E2aCwifOB9
83hYI85HFEKwLX53urCfWFxbiaI3vKVmqAk8fIl3X/5AV6yJKUcIY1F7X+Y4I83ef9fLcL+bQDzH
E9Was5U+7mxrd6tBNNqHguBvbJjOf/MIBx2+PdycS6wcQh2KEv2C1Lrf6BIEOd4/fXyRFqz6wLc9
dQh8P2KTF1TKTs3ftLXEfrVC9m2rHlOVPngMUipyvY6ZBUoO98C1UkYPfngaCURiU5DGkAJCnzfV
A0r2XbBEMhOZ6cb3B+ao1zv4apEt1q6Sw8tHqtWN5h8UBvWRRNwwiL3neZ6dett76MdOSqWXkx0U
/hFv/0WVIGxq+9I8UjvLAoqg6I+JA01+FpFGdOkZ7JKo29h+NZ/bXKLQpgypu9mTudBjiS1hjkeU
SkhhugwQ6Rb+8pgj75ghpwa8IcksXB5N3Oq0N5KjWhOp/1MLZ+Ay94wsC6tLcWDZguEr6PgEzpnG
WzROchhgAybaqID0Yb7deT9JBrkf+OFpIwFnWiHjF9vmbakPWYxYex4evx5xkn9mQVLZi4nLBOVw
vhhOElbgvLZqsIpqo9MQGjAy2zU/QOWTYhbcEIK4wopDkpu92csrb7fpAeSihsWjItijHb1LNz9+
NJFjuI1PUeuz+lO+ZubxGIaSDEF9KB7Ipz4DhmnVx4fYfC+eYJF0igW3UIZ0QMYhqvrpiwcQvZ2M
VSvJPGkr4xXyyXEbJhFHOfMbHTWm+tu1mbxV6F+DdiwWFLdc+FNHHoaF4qsfIcVMBCy2EfsUOjfS
ww5N502H1GFIvTdCNtbkU2ltN27AItrlp0FBbhvkjxTEUZcJjLlXLlXhNUgaPhUPUJ2bJm/Dx46C
4vbbcUZFLibJljI5Q6tx/+/4PC5wplKyC+35yJ8kGW+umYAdFx0T7BcfxcfOWX/qQkOIdWjpRW18
OQ4Hyh7cG5Up7/804ny4YbiGdD6um0RAUvwmLRf9TtnUqQK4GUVmzOjygSLrldJEtSSo6qV25R16
xSr9RBX6gtzNcUKCiMkW/bHUQaPDhfOf2+KnsQnzBs9D3OLUN5nvW6VqwgyetyZM7xyh8TYZKs+l
pno4XPnjTHdjcxx77+KXSKBqqGsF12yw6SE/EX1bnzCUyA+Cmzu4n4R0iFG7b1tsSRWW9Po7vFEx
fMo5tJfjsEP8v90DoVavL8ENLLsH5E9fxozbaIyTIFXYA/Bga0ka9jQdYt1DDOec8rNUqvQCRr/k
ZdAQIz6ZxtKcGVHCDziLrBWL4T7sjzJxIQBYxFwV6R7SErM043LKVSCTFJIGIupdW8QSdEWRtwfG
3BQOSr0cE/p6qr5+XzTVrTCIWeWbAAJvS/Zw86H4LMDLRL8yRbrl2W0wbrXhjgfrZwCC5VXDOTV9
R7qGMUeDz5D2ogE7UHSEQIVqqzH6QTlTxKkzInirA+lm4Qus7nS517smiMBZGYAmY6VoJHegZLGn
m+hKt1JFJlt5HWhM8WFUwppH23dItYe0nGDWtXi/+FSKGfR24txWCVgTcIXd33lp03514tPZSo9c
VLd+1tY9AB1JyLQQ7yd+zG1eeoREGKh48dC+r1sdhGhlTYTl2azlmGOI4az+UeIbIwyGgqBLePWx
+l/ldm7nLwZlzUgulyqKp9uw/X9dz9P88wPK+FtOfdjIgM/No3K5TIqid+EVaAma/T1YG9s8XdIv
GD/cI8zI9zp+xVDUSvOubfd6JjBfvsd2GCio5rsQ+bDl0AhhX6Uy+OPkYJluKYU09654j8cdZgXt
LlUSolpwxeYPkDvAVVM6Ltu8vlJGX/0DBqBzsaid8oZPt1rOFkNVRFY1swlW9iZZ1xWrAbCJ/ssG
5d9LZg0N6hx9nCvlqxrpNuD+KzvQOydkWssOF2Ks56vWwthyUGLecH6i0Gv/qsQEDVDMkL/JLTIb
IaPKczB7i7r0gRA+YoLU6qUEJotPhVB5Li6gYqjXEOQoQSlnoKzc+tsMO+aeFZhCSQfXL6JJVLc/
ooM4ysG7pBuyK3sVCWRDPmiKTbBYUizoTwqifNXM/bEgVBIYmc0IM75Fa+dp0+n3doFtZcczzTyd
nx0Y0ryqCITiRpmHNszTCgKh8ppLs5xunVdthBfIF+4MtQ7TMR8HYPEimdz+BSpHBzwqsF4lHi32
XqpwiLN0B/1lzZBxsDnkjDkXcal0RdjvXZh+CG/FMoGJ7SE9Q+fs7pPcTrfMEZ0F5Z3SJvXzFW6+
qzf3ECMf0Gj0O8yg6w60OjOsFDpMYyWtvb+Zme0CRKK5PmaaDV8j21De97eEfDNgX6ISASvslQhG
+RWxOc33sO+TKAI/HIpL+eQODDPd9uKn1jM/j2jn3DStMjRxF5QZ9BPydK7rCVkViAvSySz8Z79x
BhOp+2BMSPbs5TrLFohSmzdQ9LQwCT52zpqGxowVKqcZerQDnjVInk6WMDBAIlrK4qU0Mhd/XGl4
TJKx0FWbJD1JHJMYmd9zmTChzDsTslQT0XHkX0+z6kU+zzrVboDdvhnlZqcTPpGPE5cdp6jsQVdO
87/p5hwhp9wIB7uIy5ByKV78qV1H8PlMd3M4odbmR/sntivw6qFEOoEB9/OsK9UQ/gwHByx7oe3x
V2Zo1dryviNxO0FLTxv4j7Z21QcPj5rnnYaAmSt2NAk1cfRukhyLdNO+rAXJq7lxENVIp+D+x5UD
Ouh/GODgw36+KgNVofLcJ0lBuXhbdHEOWuhF/GkmYQQw8na+4lcDlKDvOgClII31wHyp5eBy6xM/
xRVS1ASQAfsKFQ0O8R2BCSPuVdu5yDtPRUjfSy3WAPRGVEErkt/UEcon3LYstnhKS6H8xMezBpGd
Afd59Pdl6WRiTcfXUgmBb1biMdK2P7zAjs3jcU3N42vykR9skPGbyePMtI/nx3VwaR1SDqCIGah+
g4znoTEOKW1J2oxJsbaZtfrm55svwBgf2xO3QfwOh3YuvyiJnvHGBGACfQ73aiA/3h5VT7m+KZ6Q
R1hI9wLFSoTIkYxqappP4h/Sc8rUiFxwrc+k5HDO9DrzMn0qpcZetXmw79RkgwbU3eOc3Dx2FaZx
WcxPR6g1/IWQIaheFXmNv9/sCABRP90RfuwGbjAJK8d6Gw4BVYhD4SCDRvGyLNHYWd7kRxXymlCO
1kN0d3BKg9zgFeAVrZSFFckfzlPG46Cjuoxm0r88x057GnMAlBy8e/knnck051XFo0XZdgZPZDw0
CrTLXwYkP1XCs8PpJh9OTCnJjA9Bz0a0cKfEr5mAp2/PoNPyVetHZLvYTQImSnUXe42KnRAhfbPk
edDA2dHK170GHfshLRDtxZVFdRMaf7MR6JIi7ynwQEYBDvVoLZxENBAfVk/+eSkPqBDdhzHZNpHw
xoHLPZfVzBzvag4yAEc36+kWnewW6AJmtdyQrDCT4KHaSR6TKB0Tn1I1ijkcGxInQTTYpPAq6gHM
Ux9k0sej999w8R9TfV4gLfZzqsHQDH3ZMd9pMGDA5VfD6B+eMR6nwp54mCvIwNMrbQMbKzBN2v6D
s35jgXBIix/dKVWu4MXYFRHzE0dJTgcyDcMtX4kLNmdvSMPj9JxF4flDBjo28IZ1sdcjT//Tysin
eRTgHopA0Bsu7oqLMOjRcgAG9TMioOSipfhzxY7dbZGRvgBhf498TisICUcH2ib4/N7esd7BXAz0
hn+7Fb3blzMfg005b4bl87hJwHkVYvT6b1m7xUYOUi5t06Crrpu7BxiTfZIVlJ7oNK0cSDWss7xp
HnwVlr8Dbg+KBgJV+wKkD/9Cu1pwYxM5hyUXaIycDKm9xT4ZejJspGHidg4zSOoRuSAu8NeTpxco
tL9itT2TFGzhU1NTuQ2PAiW6TFsMXqR1TcAvItBcZwT1378sSU1nhqK+Ae+Q40k0uCsvaIgxXPRi
M146M/MN3aOOBImV2oIgBDIaBzuRnMOtGEMlwTxUqlxpzwA6TEliF9VuNCmrZTzAbwX/f5CTijbj
AonEiNuCgi7I6iqsJjI+yOg8tL9+ei7yNYPHxck6B6eregug4wHPQCweK1mOAixYY0pD580LFAc7
28Kzfq1AzFhBEhSsJ+msKc6w9JHj3DavRzUtkxztz2jzEagajUViYnxG69gRUl09vC4v1r9Qd4in
nrPbbzhYF16/AVk+tqyJaDFpbXXnpN2P1QFLfvpmompepvhWCBjpG0sOpVh6GbLg/wJhr8TRKJ2/
Ei6aQYpj8Fz2Kh/zmjpF1bEVhe39d/SzLw1UibPCfRuoF5gWFNH/dxo7SRPBwkkIyw7Nf+dUCuYG
qcZtrgiwe2BEBMPunsZEshgLBt111HRjAiRgq5zKr08KTiCdrinaP0MP2EBSMUc3HLaIEsKHsvcx
OZLk/kXwWotcwwQJAM5UVxRn4D0e3fAAdXZ3ZaCt8vXFy2T3XzXRdvez0uxE0a015MK9bT4E7lJY
K+dKDhiOS4IDzF2vqfddxm0u0iY/R0iK9gcJTtMnrcZ6w21hKhhSpWdIAzT2PDOTxQew/b5+mtBr
SD6jZ7+OVgLkluG0oC5Y48lRIL7ruVRnoN7sdMHwJkJXS8ze0OITW0DOHTR35p3zFsQJaPVwP42H
zDCVsrjfu4Kj7yaMrana1hAgIsKCiIWhimajvocHP4OtKJwUHwjsu5QsjJvcOdO9zWVtNZhxQt9l
UR/qke6oHtgIFXu5j+fxi2MlbCZCClx+xGvkuaBVx64l/y4nHcViTSW1DFyGQBH3OTHUGEljDkfl
0KH4/WN7qIUfLoNEcg2CpfXya2ZIpj9swUQmT7N4mV5thnnnGeVMCsZ/IjMgnxH96ulTthg6K2of
aP4LKfv3k/6KOGavPwda4fWto/VCO/zU6TGd2uaNl9vOLFInzGA0UHtqZjEVNoWxVySK5toHocje
RBY5dohxSRPABBFSH6NRQqwdEEU5ataBOaVHMmhFVskgvAUxoZpV0WIEQyFcWOOz+Ab3GK+pA/mW
/v1oXi4weJS/jlnDSItaW13GSSUM0uSJf5dt8ICV3ILcIX3pq1GBFqtYpJUqrEBG7MxNw+Hcxks7
+KtDXQX10Xp+wygK2wbZTLbl5Rwn4V68G8w95pP3m1Goq4Kbb0fieJYCbTbV8MTTqBd8Pp1EAgfY
1M2VoXeu2NjJW9E/pIyhzqVcXGuHPFlLiUuZC0u6DDb6JzvHwDYCmT8B4t9q+xGHa9Fete01VtQH
2sSFmCq3xD96T+tlEw/KqXtTCxEjIVY7ckUnqtnfgY9Wqr0adam9gavfJUinn4lEqYtNDojAaVsO
zilIT62xMmK5ypXtuTCTJqp/XKZKtSbUBL34Me0E8l0ypKaJe74ILdzPXXqQDeWkfG6PyPh0HXQ+
a2Z93G7gwJQb2MmDMIk+YDpSeKMBVn57o8FT6on+K/J+dQCQXbwx9r/kWHxw/egoTyOfWJixRVgt
SV42mrWge16d8LsKbx/urxvO+ndxAAT9IZdiCJhyTJ6JxVnwbnDtfJS5Pe786+zpPGx2Mo4r1Ozz
lcZd0C3nWTAyh559VZYoIkDD5DlfRAspsZfecigOnEUi1maCcs24IbAR8HE4RxdXzlIMBXRY3QAG
4Dl9vzBsB0Y0Uqs+RftTjS1QO/dlFirn0Oqm5B/2JnI9Bqtc3DhIJl6Su9NVwxvho/oN1er5Hf6j
a5qvV7Vb3ze6DgVVcYIeqamVZQPaF5WEAdqMVTAWwGImBq2pD9QUSDIz241YIbBI/sWg99+3QV/E
3ds/URQlRtDTIJ8mpC7sQ2ZDjmY8dgoDKGnQfrZ5NHfA1wVJtsyy8MGSGA7BWHz1q1vUIFoTuItV
ULDpze6Zt6AaHU/52v0MncV/FBNUYQG/XGVBxApEBYYOXgVBRhtoLcO8QuMEoqsT+S6lymI97U5U
YgupcVV+kt47A9dZIJq3MGgKQgFI1qHC9QHwubfQserrDDRnGycZKJZn6VNjhJbtj1XUj1AUEiPq
3wCv80qUqANQAQtfVy/8D9Fs0L+qzw1kkcMO44OPtOKjZxADwgIAL1FZPapLM54D+uj8QO99kobj
zpHx2mno1MCbhLtSb8fIsKPPJkFjdeu3yXFE0sOWsyqB8QlyUG1LmPHKfbK7LaN+mOHTbxpfYmn/
OdIYYjow1Q1fSe0Re+pd0pN3tzr8gK0nZC2zCokR0x5TSr+2MVtqGwYixhhx2qPDDNFVjsd5pXmw
GEJaLdx9xWtZxZVzPvqh3feXbhratzDHyNQwaZHfW9J3+dYu3VZwVXZUT2jjImTSE1MCAVqe5ndj
3aNs+Fh6+DuxM3qVeIU8PzIITjAqrLhVZGLzWx9h/oU+MPOBjN1xO7K0dwLQ1NoBzreKISPMNBFs
Xl0B/pvwByXodGJtGWcNDsA5aLiT0khhLUSl6pJwdY6btvguav7FP7TJ4iAdUSC3jnk/ZosR381l
1DbA2UJop/F9xMru5jA9GApfzG/QGIJikVXrR72s7DdW56BnqO7sxc7EA5y2hl1N/i6dFzz+B0gv
CqOKsTx7++1X3ch+mZD9lIRrycgSsFOh/x9MYxyPpXeYVgawJw81GMnKCpOzHa9nctT+rt3P5VPf
Gvny/fsNLX9z6cclNQ0dH87fPTCENlmvVCCmYBuORaNz/PURQm8W7AyM9FrSEOkKKwI+mNU2EJlv
jN41mBBM5/qHDcqbKkiTYYA+pvrbbWf3/N7qmiCS+qeBfv3w+8K5kQoDAjeZAehOuQsn8daM1cGb
U20CPpN8FOrHxKjYQhUTnizVlsF05OEICW6Fvi/fwTULCEjqb2dad0KC0/ECn+MmtK/MrwXMd50N
l3PBP1c0jdwVXVJLN6mFaeakp7rClw25LWW6kwHh5J7lfoL5n1CWa0u49yBHusHhIIzpiFoWcCWG
mvhdFyzO4ffGTNcFwNWVfYIhRCzA8ChrgDyfnNfUuG4+9Ao5o+p99uM80rhrvSYD3uKKhhOHOD1r
iiIF+NlWKxashHvCLpLuTXzL2l520BaX11ZBYGvlwN6LBQqoDY80jLizAiN4rH7YPmua6h3NJjA2
FmYE7uBfFcF09tXnSowjStZIVTahOSCedg88EzolihzCA/NJYZ+onp9JlQ5aipPM4dcCNN4OPSOy
xSTpVjXQX+uCEs2YM6cQbS4Dam/eBMqNVWRnEe7zv3nPkXbMkodQ947zoO7FhosW+tEHyAmtyieA
gxHrB+LydW3APZDPkW3IPRQLlxO6DJFySeqxSMFcgYYFcce702kmLMXYrUmKf5MdHxy05JaLc16+
g3PEAVIpl0BL5gliD3xc4VpBPgWUvEfocYkwuaSnz19BgExb6nxOqrgOsk4UC0RYBPzsP+6lwdjV
LWBZadGudGfFNKAphWeqniPjmFjdkIY6HnavLVQ7cxRJ+Q5tF5MBl4n+lR2bOp1NVqDkVkywbc0E
0O3ai5YqAyqugyGEM8sSQ7TOwqHWCTuB4iZaZuiIS2SN2s2CeWrIXRMh+VjQbL7OpAW8Qfj02Kyg
eEeZtoPkyov1XapmaUFw5qzVxjDxuiLZ67eGu6Xqm6dwpBCZ6KXmYt0+nTHVf9mUT7Bw9V8fZiFT
9IV0OBRzjUJgDItItKl+qMC0YWk4+UWNSgMOgudWKKyGgOmY7DSZpCZZ7c+qoNlPVH0ih62Ic3bp
5jL4V4OqdkLx4k6IZ0Nbh13eXuhaIl2xAUHSJNIwScKgswDKhVE0rwTGfYeU9Cq0m4vrNt++Zq0g
oIxnNUwucJqiiN3bNE0Iji0MA7JPuWP5cZ2GYOaiuev6gVkSWD7zWKveP3QKROLi+xjkZP58D3Rc
bqbT8Lno26vRhoWAj8Mzsb8yqQ+O7k9gKBUKxvwrX/lrw0GQRfQIz+QYmZEDDjbpeSD8ISft+YYX
cPiwQlet1vaZGPaRMZT5sKeQCXqA00/rQ/lS8HJvZG3litBBP9sU08JJZ2nYi/ceYh/0BiAlKnW5
6vS12Mh5H2SJMhrFdUoV8O+pUNzCDmp+k9QS8YkXVPeEVzUfTeJnNKLMXrFObTf50gTctuWeTz6E
fuMdPEpV5Yv21Wg8vaqQw0hlnAaTOcezJjYLCQiw9f2XDRR++eIhFFyGEzzrEDqFTXTmmmA6N4yz
lMqG5RjcWhGVsPHUkkcEXoY+shnte16Z8B5VDh/LQXJlfLeu75V2Rb6UQVLTu05LV2Vtvp+qon7W
3VljRRKf+dX+cqfUdxMsK67RdHuMtPfFHhB4S5Xuz8ZE9HO/A6SUa0XOqGZ7nanSTKss5PuegWlR
7Q2JxHp7eI9V1ht7nacnwq5CG/tykj9hNIe33KS9yJw+7JpiKiLaKEgVpleWS+m2bxcRwVmPUmbq
F6gLaeIIlnf1bb7fmGPplByIqC/j88TTTVPuWyfewSUVBZHLGAi8TmAkgj2yL3xFdsp1mPs9s9ys
P0TNXIYw75ywj1PssBYRvfbBw1LYJwn2HycauDk1JsX37CE2D+J6Do0Uh5TeiUWet1hgKcT6tAV9
NWiBDvqs1xnW0s5aVqE3wQ7WrWDry+58VlfYtSyuWzKWrIrVuEiNxoUHp5LZ/pyff0S7WdefBvMb
am+8+U0Ccj2ZZCxPFyj7MEkTCsiJ3+5a2+exdtH0XMsJIw5z0q3cQUzS/tWSKrilUNjq0ma52EBT
DTsKK9A9OvVYSt4qAJVITGd7ctaExEw0eoIjkqJv0FhRXxQeUeydWs7mFWkbmptFstMcVqWgw2Yv
M4Gl38fiTBjTU/+Ofj/o7cVidICRrkxreuxNC+2fUaXMPSRtLF6esOc4T4M5gVZ+uB+aVcknxhu9
HLUsumwIM62BR6Lc37iV/6hurcUNa1EfCSvZqv1jciKFTXi/UMM/IChyoviA7k7AVZT/u8cLeMl+
Xxl+Rskb0Y9oqpJewqJjw1z0jeDKCfCQhqmMZzWRIBcbvuHbJhi+aU/GIv9oRyTKsWXkLa0JL0+X
s9cFg5aLVlrd4JivozihYPSuN3M0hk1seTw3WuGIetvlIGRfdYIKOO5FyU5FPNLwnF7w2AyBlXHM
PcU0pZ9Xr6Sl/kgob2MCY9rT198O3qK1tvxjP4MTnFsgYakhiQmKfZgqMZITByKPe95GJ3Wtg3yI
EVJt6V7MSyBbOCc5sJWUmTeIlz9NVUYuChP0HWuqollRfNDdTKkpvcAreW08YXrwepcCL53X7AvG
XkyvPn+HReiiKXvGVMkweksp8UmZFPER67J0ytVET67rwHNc8h7T8reG4fLrdk6A81xXrNrsdX8k
c6VU0BQ9lD+ovfWfRSpU6xR+8JgCHRwbzs2EGse8nX7FSDst+Cpk3pGsqD1JSHOeP/dtXikCSnVm
eK4RXKswBcLGPOR1VGqeJakO4oelzK4mpq5fE0FtETo6f3IpqHMmxxwZ2VYWP54eFmuw6HtDjPh5
s51sB96i5y7ftEyOmE2yXojrAkBhOwkxGJNhT1VOBnqBCiw9xd2vX7slgUuzoYcSsrKfIGmiE0ng
XXWHUKgnoswqjw1JM2EdbGuLCig+GHoIIykzjT6Yg3CgSnWEevZFIOtN+U6yI6vU7aC1oUKWTpDQ
izYd7zQb9ImJE8R+WM9r92jBTq3KATo86BPjPktYZ0nOrU1pyyjHUPfLlazh/mGOoixLq62WBNGU
BzUmhBPmxZuQw3GfPqhAAWV7xTiqHvcexaZoSjbqZLZ5dh5SjhKT/9jgVVTyBbzC+j2MQi+PIiSb
SD0PZjXUfwOlAe9nn09+Ot7RfYMlo7KzXwj3pvk40QgRei6PB1sQbz+f+0Ses1/dd78ZJuCUy2tY
Ptc86eG2Z1YOS86AnmbEMk5wzlT1gQ3NAjqsQaaCcwG5ppnYQDj8loqgC9V68qzGdZcoEiBnx/mo
R6xmUJfwZyJsCixTmwt1jzB/L+bSjP9F5u3l8GU1tvKxA80PC1d5UpHnApsBOHNodf6zreA0Vgw+
j9naM+b+2sx3meyzsmDfHB3nzCe5bqiJxr82F0yuMZN9TzO191Nf2Goom/n26/fi0DffQxRbND0Z
6U5V1u4GO9Fze+o+/gkr7EhL/CEOVpmlpLZBnEEyb5h6jRH2HqOLGmpTyt9c5XAr11AeDeSanTDz
gNFgtKpmN2Ade56Kx4S7eVMKP4U2AcRaXEnO95YigTZ36oE4udOR+mjtlfaQ4g5cTWQ5CB5vG/ts
6tYdxlayxJytMb5H04sWcg7d9jjDa6juT8DG0VWij3KRaTjggOqsstHlbxr4mBChhDXSEQmZ1PJ6
9CYcgk4F9RHeeFhvmoBKEwwABpQ2IDsxFatTqbNM+s2dq8nzVmmtzDmbh0/Pjp4aVCd5nlS5s+mb
SyOVX7uCXp96lF7IQCMVqGz6hweiqDTixS2ckRDN97N53cob0sARM5K8xV2gqlmqJhBeJvrMagO7
gNMyuPHtF9HTfHQ8WudT/bnbIhuZCxs2EqNDiB2k/wdWOUclIJSwNedRU2A2XN2ET71vX5ulOPkZ
nbxgQ8YiCE8XW4kEuOsGdR7A/lOB9NdD2hBEssCk7b/qGXgbZQV5d4qK615gQTGiSeOGPk6JcRiX
791ROmRYizeOaP5/yHd42hwKRhn/03FMKmGp7uWHJHWE2j4n+vgCL+4FvDlzrdaGun04nR2BBavu
KXCwkUWCQ02VHgm4ad7fqrEG43WztAo34irHVVkxkugrIRoFPgEAC4ZSOwA48QpUhDWjisI2Brs3
NQHx/+fmqpp6uxDQ/uKmNikjQ47T5uqfejoS1oAXOsRt5stciBRCgPLLXG3MVprbREh5I+exdJha
SvYSeMhslHpxumAC+dOutgT+ISHsPWa3CVfL+FNhQhfi8VmiBHepK6BA7xQWgqV4SOo9aYUHUk0q
KkOBghgyJF5SO1lb8QsJ8bohC/V5zwt+XFMXMXFiU/2UAjRXxD82KYAEWOdDEReHD0PlgjfeqfgI
YqZCC0YzqUGEAkCrbWP19N/J+SamV95gDicHYOqT9oCH3MmJ0/YvB8Tup/IsZDx0YTGXVqUHEDsE
AhQ6Z35aESbGkYWlgPN972d4h2f9TLYNc49LfZ4ptwR/iAQ0/TMiS/7qs/3ZZf4PuZ2QUJmNAHF5
c75L2KhggNldTDjZGIsKUoESze+Vvtg4zHP3DiH/7CG56h0K7pG9uQjXlEmK09fMgw5bN9l5+ZO/
jWBUxrFYgczPl/U7Op5Cg0jkW+gvtZefrucK/8/QqIWsX7gUUljSLp/H9Sg1hLfiKg+Ok4/UjZse
hO2p8Aiy1LtG2H5zcS7P+9jukgTyFnSg7gufp4k4/JV1P6UbYKbBunPlI0ZG939IudUPG+VAMeKb
DQcC7O+nm6hZCq6MG44TDIU2cnFbWFSt7CXlbEHEOenyZK7B19TVKVHRo906sj2dTVKUYZIL9Gs2
BOa/bfQY/BM9L4r3ExdM5VyktTKODKziTlSehDTtBBFePrwRuiSHb2u6DUsX84t/pR0RqgEsXYQZ
C4tgLO//h9E0Y/fHRtj9ZwuqmqiybJA8wXT4eo/CBiQf3dJGkgQvP/M1O0OvFuXkLZnHmdu1mhV9
K8jYKKXJ0wNVhhyarz2zHInTCHkfy03C47jCESnHiCKSg5x0iNvU3rdFhVcU/Eu+y3C12hr6lIRk
zCrq/SFW9zoa3Xg3o6oS74pw5YeEjdRa2JmgcPjjPgzDYoSaAYxfYaQO1kj1ro/rYHw3OIz+M00h
K2VvxRd/13YtDJqxra0JNmBexaAh0YB64XXyP15kRenyKXmjJtrsa07gOXQtk10l8bDw55dQECLR
o51qrYkmMH1TJGdOErQYL5pOD+Uv5MO2KfiX9FJRAOoEPL19xT3TX/L+DE7avfap/HBOJRj2bqVC
wZPYJQGeA9Ci3W9OUItyw9nNxaAeyock4mUMx4A76AT/cU2V1pKKvJvNOQ7Xzk4j2gY7L0wP+RaT
hYYDSqhZgmIAjzaEFr8nfg08s/2duRBanhxCqBcE+f01ABZt8Jf6WgI832IR7BqQKc8n6/MPSD4h
LFl46qqvx+27RgHmJnJ2I8FDpMu2gHHdq8QdOiUziY8nSogPTXVqOiznaWY6TtfphwhC1pALaKBG
v2Mf9XONr7szxPiohaLOguZKWE0ILZ0UfrKs4PaE93I1kLT1Pp71uVF+aMmurjMUGB3pOGCjAzmt
xFAeXFPy3lnav8tWICNdnZz+QahhNwvR0nLyod+DRGjOJA9r5GmHc1FRVIdU/XD1b1IRKUcTVbZ1
yHwaPneYOmThS+tlSpzY8/6rmI1PiseRJOySv6N6nsGWmei4NFjb0VjqdOUzvIbm9jIaOCI7YqkV
xQHGtWVRJDv3CMci3Lw1gBBaHiJlBuFoL63+GIMDiiR5IBVIw5dYUjmwGoE7B4y9PFmboRJQg2Gu
O1SUpE4Hb8a3KVLZGuA8WM74hQ1daI8dXFGOdpDhsEvrNTXRPQCDlJXEe9yRMC2z83JaAcrgcyLh
2Cjs5X8s5FKBBNOH5GWN27B5OjHQVUUVRLuT5WVU8C8nx1ZmSHTcBrmAH5oMT2pjHRM3i/o0mtSD
kFrQVmq4+L3AQscnXXo66UKouHYbqdrW5SRmgx1hZeFhOCTFrWt8Gh2u04W4wsgrl22RWIbUdb24
IES3lNYTxeYcTxbqSv2jLm16VAnK23R4M9/w/Di9D5B8RjaeejaADu5cNrGc48R0KI4gbTU8qnd/
yQTcsVlHBa1jNsenjMBvJU2f/MOXYLhV1lmrbmvJslmtFei9JODdPT7NpDE5AWGi2W7uosfAzyBG
2q8figQdnxAXuS0SS7xAP9KHCGxX6h03imOZsejatbaH2m4RPyybrtD1/S39oH6016ADIS37uJxD
BQKjEwiXWp4BfpTDkxPYbEvycYNQmVKX8fRqy82nolpXWzE+l0gzNqbCPZA93X4XCUpsk59Mkbnu
CBvM5GWddlt1o2s7c56NseLTW5YthjGB/XxzjI6ejrIKQBZRiMcAA2c+3GKwGhBWMmllbFtbOzmY
Qv/Qc+Cg6ZCpjdTfzveHcqWxiRaSqQEo95zHJfBXLrysCKpt02HtPSNVHqsF5iaaq3KtIhegVWU+
rVbvU/KkBuUiDLZ9S+4gScxEXbR3ffoxleqNSiSOz4vzaZKHIHPdwIWm6VOf2XNXls5vwLlDaM8u
+KxgrgIIJIcXUWjUzzE+8+2YtJU3Q3Q6kcVnkGHSLXgmLR8qv+HBORwz0p8qJqELTuWQAIdK18dZ
wTrmP/gK9cfJ32XIekz2kGSF2tKTpFV0QHktJieOIX8t1N/LfwLQ8aZYMOn7LhRl9ja5Zlbuu+z5
4hgl1eFmP8tbcwraZywJ/2YaZFScBerF2v84LzyAD/RnCbb/Yr4yGNL2pxqVB468q0LMbjpuiRwS
WWhW6jj8g3cvcG3OHPyn9aIDbVBNfmNiC0/YndfF9Ea5x+OI4Ra5+sFM87r3m3QOg88kvzFbtDR5
N2nO1yTtAbpEnMyVscMSEePVdi6Gr27ZNiLm0n5F3UEt6ZIqP7ktY+o6m8DOkmdq2NKENeq8k9D0
8BzgI8Zj6YeK773sDjS/ZJtwi7vH/ZY22KO5Ll5eqjVYDGxRjiELCL4NhJH4gnxBaSNTN6SicdXO
SIPf/3JIBJ/FekZzpPEdte/5FKypFo9iaMOX+/HB3UyWOmfwspNv7MWc2LZkiZ4VekgQmfx9QbTI
LiOjsmYSy6EUnKwn3XpOQLd6AeRq2Rx50sOC9SVRPCdeclLwTAAT7lY23ZhYciik7bdrOazyqDjT
WGsnj3ANku+LBNCaUpdLwed2GQGZMUu6/1iz2n7G/ldpD4Oka8CA9r/Xp92UU+bGBK73Nohcx6Re
4ecJQkJlC/Z3wgH1VsVeBCZj5OJTGi8uA1vi8+3khPG1E7NmTDX4w7ldYWW+L2QLwB2PFcU96d9X
hxJoAaY5FtCrxNt2HSRk+4ye0A2aQq+4APdcc+H053ucxxLrBh/a3o2v9ClNtxquC3gWwz+xasAk
mjfr95KPm43hnbGOddbHgVRW4PlSOy2V3totiq7pFkysr633tcQroKj5oWHsi2+Lak+4s2UlsXAt
z2UIhF6L4mSvXa3SvltUVS5IXaGBO373oP0tZW6i9PMwAjsS6hqqr6Ge/BadcDYSTnoXkyY//3Kk
VFc0T1E401mQ5R9ZOVD4kscC9Wryc/Q0Q8vIHB8wpjJtF5s3YpibIrzDSePxGDu/HSy5SixRHY6K
yzxzxbhiaO+xJza+Gh7rOufXJjIJSwCM9fyMto+beLojoE0ZVo3iHNxRPb3Oe/TM04judqDZSfIj
PdhXk7mAIwAJ+sTN4h7n1ac4r5mjJry626tm6WhUu7jKacExKCIN7aQGw2WWy4W60+Mu79gfoDKS
alV9bHq5/fFruMrYGv6fosCuwQQnh7qUSek5OcLbQjU5nuafWmXIjGQuKEC5g9oqUFADyj4tOi9Y
UHXsFKHCcX3I+tArfqiiXN9/75FEAT+Sb4pq/vwz5Tz0IarioQbIgrbd6TWOWTbvPGdZFBsa5irS
mx0/d6Ib3f4kXOC0zciVD3k7pmHptybL7Cf69A2rD/MLk6h9Vk7D/V3scuhB6PhEhPgj1EZc2X14
LMh7nSpz/7HLYtX6bcJq5eoV8DeV1PM6AySoCdYV/M82ICaREL1nPb/eydP7D7ReiKxnwHspgkYv
kCDrJrqJiEDtldLUjtdIH0iLrJUTobUH/XJjvcEM32yxIme7Cj9PBABS5b7UydzrA2mH8BZqtxl4
SH78D15LghGPEJJePc2llDZsU0da7NurcTsYLe/ZM43pt6tF5kONCOHeK3xN8B/JeAvnPwVAsiL8
/WoGc32/RrthVo3u1ExFm2rYvMevnVl8Lfn0/mpOQZH9eFzO9dCvCLYcPyyhKFJDs7oZzZ2ks9yQ
JQxcNlDM3WdPfcDbSd6YHKrSKcSK6MHg8zOA7PmOdTm29i+XpJQcmlnEyq7OFzK0dRfwa4xBFuaw
X+Sgz0gIy/hKIGPf9FYsDzQFaGuhwDvd4kxJn0UQp12qzRQy0Bxu9ElYv3iOPX1kh4Hf+0HOkRjM
HThQhY6AvZpxrQBYL9gAhx21lvVNJwpmpxuYIxEBEsmoIFA5bsqIGE8bwIzfdYh50X/XZQTwtLVH
IkIAwvXAOyZi9SoASeyv/LE7lF4rPy8aowYpM3SBjkbWqt3AIqhoqm60UqIt5Lp+mrihDeEhfASO
/w/WOv9JwGxybKN800UrBuEHB70tflz6aRXfn8ls26fqFM+Rx3rK/ZbOr3tdFjvuBbYROZNYwFuP
bSY8qzKGCPdK17618Af77EP+g4HV52T0cVRSHAlNF44mSO+tMVjWAl7ikUexkyyRuJ29Cg+Z4lTv
P/FZesjxngRI0/wlOI0zFXG0aH+siulArHtveRIDhUca2vS5HnC5u/kV0QVy56iyHATxB/BeQWCT
y7x8p9IuUI5G06uWrE4ySrqhZ9htC6VEbxD7W+FwxTrWV8HxD207KhbqPx/pB8F4GgzS98Ih06YD
xiwUP13Rhsvnw01VOUs237U6gcoP720Zt75L3iEWRnNBI7JRHxRV3EayNHVpBaJt2GqWPptmNjGK
Hf6Grtzx39MQAu+R6rB52u2RLB6JrXl5OqBLy6Opy12OuJWV0N2IAIVVtn6DXCL9a13J/BD9cmCN
MsIM2vUOCp8b2Atb4p79gWo1dgPVJ2c8RPG3wM6QXGanRevcU4BVyt4u7GSac1Xua8ndyIR2fe6l
/znbLm33pcl/OFYC3TBFybwfORzIhtrrmFrECmaqvi9I7JhAurwwuMRZTO7BplB5PzoPbjnl0Vr9
pVNXgD+/GYkPnRrNVHNsmDAFhx7to+X4y7iqz2n4I7wLF+1O3+BKxN01hDLrCN69l77upYrcSyrA
r5+SiT1qvEt3Zc+mH5uB+3+LVX/cl3LEDq1RK3tRTYWEsnwZcFSU3bhcz1+ZnNgRykrxxgYXBN9n
tXidiXmkMBYMKi2NNDZkEBLjLvUi3gH7wE2gbLSkVYV+cMFwrfRAx03+s2hwwmOICgZHt0da9u/9
61TWd7/pWgRD4pKGCcZIl9c8f69SG161oxW3b34PnwVdLg8WYqPItkG04oEvF45DdsU/kdTzFe8U
hSJvpYlLiTKD82HqIdCpqvEMbiIWAkijmSFDsAl+v0B5TYqlWDkbwB50vXc3lRnU28vn9R+xYH3y
ZyeANOnu4e/EL1zM1wZN6PZEgXI3zsnuBR4/Dr3AgfCIGR3yywNRY9g6SIUOXhAm/H/OaFh96yYO
+ZWrraW7/HQNCzp0+0KTfj3nTms3gpPBUd48PllzPJNzwsVcEB4GHWwa+saMjkhRxMw6K73FZ1fk
8E/mWOczHqoJ4/UCh5yHHZF+wB2jeaHruEPKqBMU5XpNmY0rIVtSle/UssFoqwI0NwiFLqJqA2Sn
NhQkWHyH4pmDFODp7JP39PdY/5UGMkr4opri6dZoe46xAW19hXS14xcyVnNnKmloprDhvJccCZFa
YTODQ/x1Tc0taD8NwMKdNC0PmFBebX0wtwX8SK/0yaWF90QI2XOBFSsIylIuuOdHaAPVdaTzjtOI
8gT1bh2H1ZT0Jt7lsKrZAMIH+4DNVKNDbkH9wqxqJcCuJLupYtVT1WwO5R7i7esSwQvXDdbKNs2a
VBeDD5RN2phSHkvLDgXsdcYVzaXM44+bmMtUcUwlsDgS53+88hSzUAx4ZrEPm0rTtSDa6pU5bMgp
Bg4g2ZT1OSpUdXhLIxW1G5k5JQ2htG6/tnUMgGBmxBB/awsCdwgq/UIo8ejV9Pq9D9f0rM2nSNAG
EOZDjXjsZNclIbyv/ZjrAPVYuk7fvFtr/IF0IuIxw4ilPGof7xQI8iH5CsSNFNzEoFApIFQ5++mQ
wkh5Ot3MUmOIdWoOvxfWy0kZvzjW2JxzmpQNqDuKKzNL0R2hzmKNVJHhHYHeB9B/11Yed4nbCw7N
+qlhbIIl+POQwnjh7/cHJN2ZeEI8B/TcmHsNXdHU3RpeQt36L0LR7KS5kJEgxe9MH/NYc6oA/1EX
T/ytyN13h03lDvfNDpHNLPZ6n2+TAGByxWcvRMLpMbVDzI6y5gXhiXV8SstW5TwTMyQ8LLo8ZqgP
diJrZnYt6I6mriJpIRN6p8BG0LPgJoCp2LR+etlOzBxQCeS2sFsgWLuesWO19gfsBn1pJNX6ylQ1
4IxA/hhpaOP6rlXXEynTVtAU+KEjD5AgvCyekRC71Bt6DIlDsniLf1AYGJ948anz2kQOMtbhd9ey
M8vmpT+txNBoe6/xgHSvDpNxRjw2LjvvSNUJPy6ZjX5Xx7HLGLHqKsZSEtd8D6+JcxxqQJ4FVuIX
p2U/XvcCo48F5XxKEO/F1642CA6eHjC2sp2oyXOW4nZKlRMPO29hennZNe3abtMGg8t2GnFa60ej
57xU+eMEdaIG/tM0KRcIHJdW6JVITYi0gwAfsHPZQEuFpg5tkmUpHqRJMgp6NI8MOzUGF/vHkVo6
3vtNmlE4gEApDEJJdHpDJB6At1nVr4kSdlBONO1KuH4PJ9pI1Dy1tD6r/XNzjx/P9Q5CtZOBcvnh
QKhVFRrz7d3iitCgfBTx+1kg7lRMYaEwu+SXKTD6BxzGGzuOk1TuE29RY3tLwwZ/TVSZ8BzVJDIT
DrOWSzMAnma/6GztPXeI7KgDrzkrnwEyx5BerpqEN8/vLm4A5zSYB4RtAAgJHCs5c5FhLQY3GlFb
RmVhGShKVGvLrrzX25n2wyaaGMm7RL0YtchmIpHkj0X/OfYv4uOImsbmWPAkZwSb4kIYQrqLmInY
ghJToTNhM/W3jT8wGuaz8liIWZrupofdeelYUxytq8l70nqOLKAGpiA/CaMHTUKnoRbNwazfpR53
JDNJ/t1FRVh/JMOyBZVPIT3dSwum8jHavNq6cUb2CjbjGjC7wwsO7hkZQe24vqPn1hLbP4Fo+Tlc
kCGN8d60LJzwHNxe9L734yFi6qVXhroPCezwkEunY0HdKLyceCaKbVYCI9LRefNPk2AWE5Qss9vN
KxNrg2hlXTLXZi0EetgJGKyik/wEimk1Vsj5dQC7eTAHjw1CBOIRCbG08HnaljJ8Tf9RBGLjw/m6
FPyjqJRt6mJfo5GdTQ9QrmgAEqCdoyW5TEQ9DilvSLOV4SA02Qab17gDRP/uB1YCSuuxOJFigYMu
JoOyeOnmtgG7i9hsfT4Tm57lCkuBaWBhVLyk4hkTCMZ7udvLiL4ygGMDKamNdNGRBicfIeg/CpUj
1mlKSNWhS9zxI9pvIGuaGljfvE3Jo4nmrCPFX6NxB7vNCOVGcChKyS7I9G1EsauZvPLsfGtW3yDM
yEAmCpBxTE+XOnGn7+VXHhr2qX51rjAF/xZnym0KmHLcPQu3x1s3Ut3TWcCrR+WJ1cNJrCwdDKWt
jCo7x3B3aHFQwKdnRKXHKuk9etqcfFnVNbh4oiqhhbX+4RrM4rdnzn/TZQ0GE1ASGY5WhbsrOpmL
yLnQyA1+8lb/ks9j837fQvmfgmcjB2pZtRRU+VmZmrtofYgSg/nHxjQj6V7sxfw8tH3/UzlxrAma
zG6vTPRmE9zpIQSwrhbVvcO3h2frYnkMEEZaRcY9UzH8jlWC4UWV+VFSM3Wb6B8OHioduGIJBYpj
Nr/+eolb+lzCtGhpEO5MCtKxSUQEcqATogd44yWhaq9YaJ2vcAtTx0W9U3vpNl+Imf4FZo//+qyp
zpEwqqqEm16YyNXxuTveYwPHO1inEPlgUt122YokDLjmGElUBcurqS9Nq9egqdJNGFcJhtnxUrXQ
HvGPvqjw5lbNnpfqZCxkAscU/A4JenvRsFj4sSMnueVnVa97HGpnSjWBfxGCj+vDJAxIyppcRqYN
NtVQ5rFz+7DI+P/Qe9u6jnZmRG7rxG1FCEVuERt8x30mR0U0GVcR+CXdAsYK1mpZfMY/YiyCyASS
GsVCZDnd6RaLNpVxPv5wKWV+ZmOb7vw9+j9kn8RwE+4cpYfIKE7jSwLcEDAKqPubKPf06AAWdi7p
tKQLGY1kXCBlbzzb39Tc+r6UYCOqVryNbbBO09LOnGjwEQk10c2cFvw/SAEz5MU84RN4hDkPFhUG
SKullkadMoCWNlJUXuXxUCpU1i6iBvHkb42QSeUIXSOVGzdw0gDH0PfvKXdCfHt2pPdkKkXlsNuq
kB6Cq/zCqdr/8qZEqygo80pLOm0YswS5AX7uhwVEEP5294vjGqY9UQtEYQFUbDjWOEvU11KqSEjZ
i/56uM3jznhrwE0fwtaxLNt/aAO57VSR4FGD8vR35yUd5Gun5IA86zL0saZvIfzt+W+TMY7XBZmj
9mtNR4AX6Fz0BZP3kNyFbtlZwWf6zZtbR1EyqvYIHwCaLV6xy3FeZsL3wHN59tfTfjyj7aSFWVLe
WCVM0rhhnyvlcUjK9UeY5eSLnA4f0MJDdlbzMDGnm9QT4AqgEIUJISceWKjeIHfFCBA14th+h8W+
XhQqdc+eTpLRroDIFWxEuZgNp13XpI67KHaS0njnUqHMxMhHPj6XqXW2he8dP2FOeTLlr08PFprP
5v8BpxovuBEcxmmH/VLrudgLHvwVQ3lv++JE/h0IStXl7Xca91BXAe48+VwGI9MiScDTnw7gGV5b
kZvPF278DxzOHQPY/Y0TC3QqzTkbtbDb0XqYL21R9CkP07YVu3aPrGsDJ+zOhK4++P+I2cfRAf5h
BhDKimP6QcrPMTzzLhVpceCfE/eiYC873DKSEkygG9yDM2H9Z9b39b4cHQe5uchJtnkA810By/ei
gh7fTVHXnAKKcsfoCUvkb4pgBwBiemD0V2tHqzpUQxIbuKbtDey0X2oblVZadl5XhvPSOxFCC+SZ
2LwFB3WESXpeqTWgMP73gCnrtrHdpB3/wveaBSLEci10fNx5RXKExD8dhova22jMum75tXrd0tqq
bzW0n6GKD78cs9qQdDk0OdCOkuqAiUe6mbnXvuZmO0vf9tZoKZ5VMOuTXeAtHxgBYSaw2gNtKShP
8sl8VrMmEcq98fhdTqPvKJ4pddwBfECkGsJxV7h36jK3ht4hdD4iGVszUugfNGRvKC1ZyXroWi68
xyGSjeFxumlO9QbHXUtZJtQ3SAZqCBfK7d7O82l5L9QfluOieNwbhbn1hKxS33TOi4txOY1ps1sp
t55KA6OqeaVBke/5H4ya6aBilBnBpBzeeulivWWW2DRBGbwpiQFaPwd6P2vRHwfxksZ0gWLeXVSu
EQRPSvyENWsAcoWk9aCOlc3G/NTNuUDSkWh7Ab20Pb/CEozb2ok6Lm7nounSiW1Js082MnTtYfX8
NCa8d4dB62tzSgJNX7YzMKSGhjHTRXj99+q+HvT3XR4idUnzIeRKJW2f/6ClXH4Kl7kqQJSVe5Nh
olSQWl3RASwsyVaMFTkujUw9TSA9r/jsS6PhqKEjFMAmWsOOmMA6oUdeZlrV0BOrjipjGOovHIez
kDSjFmxdx3ck23dCfl1XxE910vkm0PCgmBd3dV9dy3w1wywCVFXBzWVrs5MUrK1tYndLJjtnOqpS
z7l3TQGdL6YhDsFUOlaUGT+uuZripcr/X9PexdCoNobvhLqJei00Y/qmZc+TNavUtpa/x7r96OD1
zW4Qkk17tW25YrulSDf8k/bV32zQKBev0yYJk0E+uyFoKc4u2mVMFRyX2rs/yhjyiQB5uYQSny+Z
hfT0UGdYL7fO+AVr/e9/9c7Bc8+T+aAoBIOLzaLRkeYwThBazFOYVSFyU3qniLf8hfDqULs5xstb
L/Nq/nWutWvh5+S0vZSH9kaC3uZIQSNWmQxpHviVzXQGxU9lFVroBXFq7AwBAZTgvcS/tIZ3WycE
L1kcpROoDNXQ3WocqKA2tEWnJE6QBHtztBlUegltnMjxIkoTrrH8jYd8uY0JP25rx1Roun/rJzDc
jmntGihYfxLC7UD6SXYp7H3MDtjU4JENlMmroeSNXP3V8v0OQqheOr4BK4eck7CqRK+4sCU4H0ku
s+tGb0Yz6hR6tmEWEIc86Ejp3Y93YgcJbKTBPvS6256pJeqj0bX1FZyz+czwpl7r3bwSMgt2g5pM
Z9M84+/vrE5PUAuE8fOj3AOjiFemmaQJ9GpkVERE+coog4jIUnkJ6TFTOHKy/mOJhv6Pn+V0FLFb
d0sN2HihLnX8LoIxPJeDPqhRJ8AY2j52stLRmYgBcpkqpY37zfoxoKVG1aWTABHeV8rPBBe9e5v5
Fv6w8Sm8qAJfetFBq/4K6GOrUtIghnX3sT9aJHc/YNt/RgkYintYY1kbdesbkrkSgyzCRx8CtDu+
4ekdVP4FKN+5jup+FfSQWlbht0jeLFruhyneeXz+12ovnP9DSX42zqWoVYyIP9sgw9FlC12/UX+X
Uc1Qtz5CzhT5DNR0tJtzC6JaTaDSJvJ2qzBcGbWVZwDQxOJrcgKmtLasCXYEbIliQBPjD4Vsyfn2
sgpuWyEN75SKjYFZHjRaJ62eL3wYW3a/63f251kdWbqV+OA7dqTzLtrIcfRtay2jFDbQqA7lVWQ3
EWsyMZQQrhZUjC6QwN3nV39FH7k/nLzGvaYf4zLHubLK0OmICeFbbF4mBQWGJK/GhwEtuq3LAwTf
yfm2EMUOa19OolB8P2ATRCGzyKnBoAqVOWHtaMRMHzxOrcEtSMacUxt+e5Ha4IwCCZySQWagbr7/
aZwGjrPwTOTp7b2MLGfp0nz+yW0PokN+gtX6IlupL+6CW1loi99ID3Mj24YjAI0znqz4KAxNQnIi
TbaAkgN+NIUwsJ92xCJUJTYDoRfnx+oTaI/tLMF9D3W5ddQhvN1qrh29jkyoxDgHNpZxBbla61qW
DNz6kw0VJg4u9lF/6Umju53pGHKEVG1CmK4lMlBQt7j82vJlAGAjOc2d1wOqAzADqUspnrAb7mac
PGM9sefs8AbPwXhIyIHHvFl7mV2rubVonnseHvi7zqxYg9UG3zShXthrtq/cYhytjclwktHkwKj6
io/Jmv2y3jNC14wcVbuEM48ugnr7ac7F6/UGKYntiYIJEzC/aUNc0foCLhCKzf1IK4ZaNN+9dnxR
k+LCKDnFVNdIYZFpCgj62ZKObTX+ODY7d7hkgqRDI1wxs+c440MwaPP8yktHm1Vmmq1JiAIrtw+e
WWxQ75g0KBE16yLNO8SXZ2QHJ8uUtAYIkX9WGncbPmmF0XSRNs9TEUEHagmEMUpSVdAr7GBVlyrz
wAFOa5rxJTTLIAnNIMsR7FMHM4dw006gdFyJfUKv05O1DZvJJzAI87COgU3goUO8NF0TKhv1kv2x
J5dk/Zu/thtMVd0goEZvmZdSB5OKx6sry2zYia/njDOurwSuELmXvWFMWzH17gTNwuayo4H44CN4
cECYmcU0t7oFRidfk9HJztDtJrrZRdbd0wVm+PnltQHSKIHATstYhfSUAnsklGRIBvBKeEXmVxxJ
Xug9Is/f3h9DvRiW5tz28cF833ROjHVsXtNaB/bHGU3BqH5VHcoGJqFnyM+hhLCZs6sKSSREVHCW
7ncPosc0y0/flYnC5y2y5pXHdVIR+LZeEjr2yaFJXFJr+kf0eXn7RgxVgNfLz26oLaiOuAWIjhu2
ssCrWviQW8T57IJtZzQXKE6iMa9ZIyv2JphKgVM3+6zQ4vMYj1e56mxR93nYendvjnk87Wrg+P0C
wD+Nz9Qj5xfQ9FxNlXi9TPQQtZgMHb4KJhqHzpD/uUKkjukg1G1ftCtNgw8Bq6u0yKbo2Lmjw67i
2yGgNprXtfLAEOmi56WyELCqVYNaARSpkbj4n9/Tdpe2yqnKmqumuswEcv+oDfFZAqg/wVCGrie5
hhtS2eLSwgQNShmAbND7rT/2F1p4wW8o0y53DQONPSvFn20lB3dUyv6WYNtb3x2TWi/+B2SXOMIm
vSxIjoY8CLr3n5PODFcr4/z/6LDdB9tCorYIRJmlPOsQIv4JrnXfhVqWWMseussOqz9XwJKO7VOY
PXTdgeZNjVLLR21b4pS8YFd/OGPxbLd3+cGH4XaniF0F/K7lmKa1xt7j2vNCbMjtiXxIfEtrYGwH
HLXFmUZ2KaM+UKazcNtCVvlyf3nwQlZi2lKYHiu8kgNhSXq3NQVDLU0H5HJonapMJtlygXWeCi97
PM0ISIRjyRuUo1aU7XHhyQ/209B093HYVRTqBTUBwmaSaQ3o1VW/yCQ67CpZcu4+P79uv9KgV8kL
nzTt9lgzkJeyqKL7akWQtO7adpv1snlgiq82N9h1oalyxu2RMyErq6g3EW/l1vkhMpB+PACkniWF
JuWHbKupW3nXjOaHRZWnkg67Z23RleUBfY8z2F4HiYDYedIaKVP4Zjer8QrcbXVXW//XkE0lZQTA
0/HDQtmq92l1fXYfAw3wcN47xrmI0idzt2vsKQt4ifEnfp7HKJTahoJjopELiO1UPItgKsJjROf3
HQHjCmUjy+/5TU7r0bsOJoLlQB+SPRlzcQ1qbZQQE+dR2rStNNw8tW82EzsDvWGlnbUE0NM+tYvg
myVf61c0Aa+FSmwvPN5pOrrhVOBJS+xueusf21aYQujd+Z+9jf5gWtVVH9AuVFvrc7jhM/hpFivM
50yShCq+ClxELUwiq0SEUAChYjW8IvsoFsZuDfkWFUSRUFWRuH8GlGstCwHzcWOsIXUga51U2Py8
x+/N/H5D9ltJmRbp1awtzbSBWP3BdAJr79rOwqn3ZDUStxj3Ut68TcJj9puD+0aRYg456gCQ8xc/
B5CtRG3sORwGm6pYq9Ck8N9siMZzDnnkqUovwPTsW4UhTQgZ3HqZ55lI1KQFs6JjDQ0xDYXdQHM3
NT0L3f+ptkFrwUkSyUXZMccAxVy/01tdh/rZ9nRfEWiYEckXcB8sEPV+YhyktGboUAmfZBJycGuw
TsomO5oTUkkbzlFJw25gIOQ8FbIYc1v1Tpde7kOFJwTCDBaVUsrGCn9STc1i8s2cJWr+adKmK8XT
KTKmEBlNfZ6o7WzqBu+fuqjFZNVVUuGXOMr5CWFSosBFXa6nQtnqGvb2P3DRmp6ef1R7/pgIicpo
PCnfNGpBp/ndhWZY++cGaYKijzQslq0gSME21MDFBmnHjy32PLnaX6wQT+K38iWFBgznk4l372J4
h8bBeZI37c3RQus8OBiT5kivqzQlgnbcW7hcT0ibIpmSot6ImzLs8U3/yhT1uTxgvUiqsxCiHaYN
OhN6ndQ/cBaVpPw/lAE0gH8ju6T2n7bJ2SzDx8fpVuYx1IIHBbSOKYRmIuDGcDVd98uxDkfigmJr
8AHOf/F2pJzNa7hw0Y/e1GIoaJbdZ/Qbfy6jQjxwyFpE+8p4GRZIj2zsMWM9IKDVv1N8QGkZtbs7
ZyJwKH8ATREIKWDeHi7NTVflJqnK9ffqyDKDZnpCqmsXIbOXV90zS6Z4617BE5mGAtuCfaNfWNSz
5gXo5FuUMcBbdnjkggbrI+GWMp0Sk/RYQvcMrwB0qpwIFOnrWm58jENSv2qgFCYPrMP1qrA7nCFX
/jbuukKqoqqIUo55+hxoNxa3VBj0GT2X9KdbZt7cjeTWbCQxYu8Q16rLj2rlSFbDQ/kF3jd+t5H4
MGBPcDF7JsiuNLVqiJG8scMD1kz9dwm5wGdEp+LKEs+XvKE/UaT451SRLRO36mSdLrca7a27nHqP
tZQRI+A9nqsRVTD5hrrcmUl65RrcaiIedRaucunZmkM/YVwk0i4+OeOEKCpqyAGri2L9ohmMWnz9
62rANemyFMA4HdB+kAKUwJFW6k6676QVG5zqopsH9dmUbepH9sZZPzsXOtPF2gQV0r0qsD1sn1XV
u5UgNYQJodYomgFanVCVQQ4XYxcdKmw/nU5vLUnJYG9zaGsP1o6jsjEH5+MwhhQPuu1j74rQvlyJ
dVyOvXFXvNUKoY8HBoI2vEkUdEULzzA7O7HaS5kktyPRDksuaeEIzVyS0KFRuO5yzp8qpl88tpq5
Z469oTkfuDVM8Hgwk9vn2QnUS7wCHX1RN5H2UoCvIEoIqFN3wA1pzbXNihvPYmWpqgvUd7jlv8lA
pHdZlP2T4Wvl035jk02/ThmxPFAF5jyXbWXO1rTEWr2/OMHBYdDnZlg3urMnAlbvPmagQLNO2/aA
uMpEdVswiGoLZ7zEiVcZjxgoxuKvKBzeOuEs1T2sNH72HZTHfgcuVal2WrYM+RNgdg5kAENMX4yT
AjoHoPDu/Gjm6BNPmmcUicT66uCm275xouq5ai6fJ6b5coyixWidMnXDZrjZicuYuRtiZgT0fJOY
1EWu+IcYrVTIo/dF6Vm4uNgf2IS1ASWjsf98dz8RQZxaxFr9zP+GdmzPwrk4mtZC88EQons7A/D7
39xPK2j1Fom8OZe+6eCefML/+2B4/UximoexfXwq/W+TZp0QAcuXv3m+dIie82VWVgU58I39iYon
rgldqoHJU4AdDeH9LK2J/mypYVsVCcWxGtiJOcX5JtuQcHwFYxI6z5a0i+T5Yzr5NkZwrN2F6Ah2
Xa6td+iObE5UqZsCfSfSJahqt8eoLIoUCcXJ1Y81DV466K0Wdj6zfkDBa7R7J+AKQiW8TXSpRtS9
nsLgwL2zZjVcLgBBhhEJvNWb3tXlsK6tl0qFb9jA4K9JwlqwH0tXYu4LMz6PD4ZEGxMbKuDwPz9A
C22O9I3n/9EpK4tniCK/kG9atNLRKpLO/Gx5PVFoQdt4e6YmmIldyppd203vDkKcUAPI0xFeHtvM
qD3qx4EKxpQEJ/3U/7d6J4Kll6JK7yoMRDdzWlkzn2e1n9rT1yXrcX2TnkPAd+3R/3lhJjStFLUM
/z+KUdEiM3bemaUseopQGbxW/SsDmB96rqCawyZMjCswFgt/ABY26+kSopPOewnrqwi6DWbOQuwa
waOrPuPQr9Ttcajj4YQBkuLEMky52oakk34eURFt1qmWmtyYmdvPQrxDWCgIHh9rb/2Dfmt78u42
FbI0xzZTTyLAHT6AMBBcqS3WqzwFsuHlBGSh5ziWt/vaiTzljRF0EYlyA+OFas+W9/aNETZ3Kx1v
zlVBTixX/SPLRMpm21mvXdMGDd3G4YQRr5vltHFmsDkR9MH/v56HPPA035p/RKTZHL3bh1SkuxY1
FyxhzxEssI/7xlcOfEru/cbPd78rNb5fCanqGjuMv5TlozvIO0mVgYVbwmSHzycQSg4FtckNC/e3
wLTqgctneJs0JLtEyXrVqZVoyfTFKFrvKS2aXStGNpl3E3y76RQ0T/EH0LRXfs5o95ESNyTL5uDU
/mJmJnZbzzQhR44iSVL/iKRpDOY3DRatCm8GmwAX8ktDdpLiEfYyqerR+cS1yEXXvmT4aF5gFpBe
984++mTdqSKV8bCX2w9hw99/j7sd8OI+Dibhv+YHegeBVb9h8h+AhcrfNRX410QRYAsfr+JiW+Zy
C9NvUFpQIRhv3hvSCKE/TVsBdB6dP5+tor46bOEA0shRng8xIYLlv2RQJh0n+uE5+t/pyimrokdF
PETJsPowwe9fothiamtJhvPWGt/qx2Yut1IS0ciiei5ehnMnyZstcmJYzm/X8V/hMjIr1ViyGg89
bPAGDSBFsFp+PeQ22/NO2B4k9c7utVU15mxdbDCosH2R6rDLeoOeO9CUUlSMmGCoBGyoJH5IUGqV
Fpee0qsjcMnRRfCuS819T3oOl9sHMzEbTbNf1+A+2257n0mjSPFgy8Olr2M+wIZRAR0jq49JlUcb
NRcRG3DXgMz63MzwUdBDb47npM38l9/I9gso/5aCQUqpMenVqit+8WlvojxcwXA3axyzInET/BWJ
dJ2+40uPGyJt5O5VI7cMxP6dtFhz6SJzCNMYXekXnLDURHIA/8ohOFiW3+cB3gVJw9tM7eymLdgu
VPb4OccWmsIVRALtNskOE7XC8U6j5huk5nj9mbeQcEastAzFOcT28n41fBprOZN+/6M8RQEDpE45
giJSEliL/AGWi9hlWwpVjVNm6idKapVK2y5IJ00otDX68Ojne0fq51offfxUiW50bpXfs439T82D
FBjGbFnWrl5iW63FYDhHiHcMNwB8cWG2pq3iPvVNeLcTmWy0KoQtwQyTXuQWuxB48xPq+2nwNAPX
VdST12W5v4ZVW+z7KYJDxWNBz348M5U8Qxbom8V5oXniOY/jYdEVHnbsqhsqx7ezZZRCiuQbuMHs
OBUZATMbaJCVbJ0qZwirhwJoEwvExiTaYCzGtyw9vFTjFK33qPq5Cyp3xlkT6D1+u8oqV3ZWaObT
Ue9Me8zEzX2c/RTM6Psvd2u8HtT53e88U72SxA0yY59o7vENdMIcoIFucgrxkWdNeK/3BmnjTV9R
97T/MJyEI5Vk6o1LLAK6oKkCNwM0hN4dk1az6+kVUNQG14bX4Io2nFcvWKrBP7M88jffzxk/ohUR
xfyyUcZK5IkH50vrBG2TNv5RXjSS2XQ5ZoPCUJzzi2573x968SXd9i7WxSWowET5SQ0tkX1YKznR
TDkrZD9LY/n3hfHOjnyLWpqz/gf8oEz+MRgeJbaumuxNJMlL7eAMsvD7KSVbfw/2ISbef+OS7VYr
PaXRx0j3wb08c3FEEFnm78te68UxP9zONstX00Cou3nR/tvbPU0wP2ojTUdCkkC/nKRuGU1Ofij9
C4uI/TQeOmclq783TXUi1jep6Ysy2wMtK+b66BtllvhazPX/kkbbzF98Qks6jSTsElxKWzGjJyns
qqo2kv8ftYam736GGQO5NDXy4kn0o8gxre1laPzdRzESJZucm+fOXYktGrQNbxZ+JNPlJbj5Yfvr
gXr7ZAZ53sPlHvjOV1ifIMwMlLaX/Ssdf2zzhJjJmQLXGpzwS3K9h+iWMD4AtFGMxqnM+06HAHnG
qndQ79hTFwxMwXA7/gtGOeMol+ooqZ/HbLRha5C8RlCue32o9lR+aDuEe9sUYgJ/osani6zpZRBu
164smvvugkimYS2DkGo9XNibGJLcokFZHfsTRcZHbhKfB95hWsP9onrMAjr1dJjkyfT1//pNWNln
exJTofFfXHkCs2cSZhsCfNBg1iQ0bReOWZzoF2MEYr7OXoMLNb+VUP6pfFzC/RBirFXrNNnh+X5Y
/qOvrK2OGdw3FJx3AORA1R7RG6s8JadWUBKSEA7pYWoTFZWNEjo5SAS36zJKQf+GPxJCzvK+SRoV
IxCjOGSmJv6c8BLS/FDq4+PIXrVJHcyCxLdYHWvDmF+gAFzzgj+ntWONh3cyCUc5lNE9i4Y9pavg
by6mRcKRktGkilZEn8CG2xh+88Un3cQnF86PLLEl/N9Sj2xiWKXuZ8NkrBxpXfjIYN26aU/GyBTm
cPECKO5BihN8oMpproOMJhQoS1yxdKqdxJPbwbltPSb2+P+CFyTsImYjlpIZZtIIayPLXxg4lTX4
OtIONWnBh0YKgz6CFSVweVwHckoEfv41o1OO/wzJqeE5fvy1ODOLFLBedjVn0Ro5oslb1C/yoImo
+obV/2jHvtQkE+cQ5jFYT/0ps1lbtEoxeIrg5N6eg4DeJsjyGHHL6OkaR+cAlAvj3kDeNVPXjXoI
yi5twwcY0S8UOwkfUiO4/I8S0+jzLXL8eSGbiC4nJZa2+wKFZVR57DJL+889BfPYZvpQcEUgptpZ
4ke6n7Z4Ajec23w5viuvn/XwLh7EgqsKby1JuxkmiBAB31g0GSc94eAcGBf4ewEghWZwAJ0VQbr3
Ke5+VaHjq+8/AcBwBQ0hCvraohMW7nABvCiEGXm5vqSlCv2ZUpbciogrAm6qvosig6HppEGXd1R2
lioARAlE6ZrBjpWoc46RIVZ0VDOTqVr7beG7wGHQ6uwG9Q2hNQhfydjwbUxXRt2lWbFShD5cmzTS
MdA4AYnvYXh8X3Ww1Vc0ISKnPRTZhsRNHGDvasGklvQm24NeRHMrqx62UkPm2ehNnxu6rpdkEz3Z
QIRwtFS3vw3RlXcAq2ZCvi2N5Uw89HlFNn3qWCsRXFjVPMXtx2/y4MswhDtbrNY9B3DaEJ/ecdYB
tUIjnHgCBqOvl0JILiU5MJZuljnaXgyrPgRTbq7CVQJWh4wCsijt6T1a2pQ5XSP0rbxnUYkeyeQ5
SuaiqUaE1s2QAN/D997moT6h3TlBVxw8xDXkUNqJv3Y6fwrRWwzICElhygMdW28S/9Am5ZDMavGT
7EYb2IM156DglEyIZS53TooWflULc+gcAgULz3VTatu466/CUjOGsDucco+xv0SodQDekyU47u35
OspMRxBa93l5wmbHtakDAmO/JL3v6/0y1Rw5oCPpFLBoP8lq9+pyF6+tAohbwrHYbi79sKbCCukr
HvHdkj6lN/bXMIRex3xxasM3u6/JPi1b8rdTt/fprAJrKAisqtVpcN9aNlDy5bxFPew4LzHBvssM
PFSbeD/Ch40IxBlv6KreGoe9UEKz2xZXb2kSJL1DkLSWxoTyIwtgwWHOljQPa/pQDLop+NhCVI3c
8fF7LhRREStFnRC6aUHZr6LcuyNwdAv7Msw88M8QRkW7m/VhbSs2B50Zf8j9en2avkW4Dj9X4eo6
GXejKiVOUg6L/IpUy4aEfcPELaUzKL6c+qz8DhRjId4Rs/zhcc3mfYRRXTVlmHADVxGy4Sdgt41J
Qb+zALoCT6LfbzKVm9strFk5+K/S+d6mtGMJGRpaGb86oe3Ib7b+Sq7lPVjWNipathNO9fwV+CiP
pS0MXKFBXRbT4d2MsgyWkS1KsynCJa3A9jAAPTdYcWtUbqvIKaXkLdQBx5f8MsPjAyB+/3atefBh
SN6m39faedT0Hez3ozM6rd6fH9gEpAL+uziFjcIING6f/as8bSGXWcn5kZBf9nHlqqJN+Ge459cC
LbifEiKxtcYL+a/tdZJHl3/xxVpBCZsQ4ZqFH4E8LHgTbAuutPcNlnBlZFbCH41aYyst4merg778
pivU9ANrefPWXLybmwHB3ycwRyH2009VIu1LzuoeNCx4sDOcPRCz4Sf1xinMMDERH6de54DoZqY4
DwJbqOnqONmO5kdp9ZV0wlMePupq3B1WCWaCRP+Qn9S2jr0us5MdJaS2sGWhaX2zlhLTzahYsEfp
1CS++E8FWXTWX4yswMFOuTs4SuMAX0i0ObnOBjaYjrL1mhju7PQetXR9kk0n9lVRsScvxHpoVbeD
ZVbRlM4pTF/LVyELTxEBzIy6p7AejDEP00IE6ZUmuemV0ggHedivlM498XBbMDg4EAFu3Jf+T7il
ZJjtepCJyjmK5fePlfh21wzBqqIfHod+7wQNezgHwWCq+/Th/MCWin+4jQzq/UkL+LVb1Kyk9CBc
pnc4gBr0t9EnA/T3i1fKlO+XPF+wrKUWUgfsLiy1qqq9p6nkVvt/nqIWQF2ohZ+eU+WQRxyRfjRH
x4862hDYHfPyHimAu0El9Yv/iBuOWAXCkQk2k/D0rR4cbUg51VIlbLB95nv60C8qP7gDrLKsKoXB
fbfA2FxWpwpIiuiyWO9g2HwhNOXt5UsMQsWMdNIspJhTs9ahWf5tRSmqlZU1pBdPFs7YOw7Fwn7O
oVJK3dc6wSa+vc51vC5x96kuChN6QGYYUf2QWrGK0pdTgzQyl9MlG+dB2M93u9M/IoWMMsD/qAL4
jQsxaCUU5xAEphikZnFJAeT3cTTcW17iBIZYoUXB9DSPddXbcFUenAxfstvA3jfkRMLBjbbjN5Dl
y34jN5uTAvgHtZIFfoV3P6ZNwxrABRZR7BDH1BgrMSE+r6u6fQ8YeKmgxgmYr5WWFXVee3xrEYa0
6f1lWNlratQgirtVq7/HVyOcJkINITF6hwzOmOi+bVc5fNFQh1X8+u/TNtHANjrxrEaUzq55JiGg
QyWMyWd6bz8mcXnL7QhbqCAKtVYFeVZEz0SVVZfekomuyBcOx2yERvuvohga6hnjf9GjKGKtD+DV
L6hnJCYfyDRd6CKzvHtPXSAwSfyQNmP8ZG8utWHpQiWGwJocfee5J7eAmbS0nEBIs4jQXfCwr24v
p3LZTTn+1TshttpYlwfxwzXEDXgme7lyD3cNpEuwOHmC4BBFV4rN2SCsmmupLa75kSG/3GRJjKgU
sT7xYUNEBYskZ++bnPb+qjcLOYpVUkvX0N44f/R2hW7LVDhWbuXeKRSRlqnjSP4bEygcG/5UcUAN
G+fhlniBMprAUCmHb2VhRwlC/xOdacLD41SfKq25M3IKdPIkrCN3QI17tDA0LrJpULi/SKZeSPjC
AwnD2M8csFGqOWepXM9W8VmOObMeEYL8RrjfugO/JhCXcz9nW5T6YVsLt9DEzqqQMVg7bQIxOpC6
gCyL6uQnbkHov3DFLeNXM9JxIpUqYhzoHm28pfmSjodvtOUE2TikCPdaQHgKXEwzpyQVqcuKEwbE
pKQvYHUsiWG85IhOUAHDJm32bDgFe8u4o/ewGJunf9XdTrhj6/bhqjANG9bdMNf/Dgad/p0pHk4R
4CsVcQ+N67N3ptKfxzOhPU4YL79RwRVhVFXRvxFnE+uZPkaBVIgAyfCncNvexh8c+g/+MbfVpQLj
iF30gOk7U3qRfa2vbBE9ZaJsM9waNI1wvAYD/m7fH6uDh6XozKtw+EMNJocc7brNsG4SMxEgEVT3
kNoccbasueXxNuq6NekVswpJPVivn8a53ZaWQHX5vbZ0cQCG3PgN+RSZcipSIuWODKPIDW3aZ78s
0vcEexTFkGlc7FY4DEY2kJruraIxkVlMbV8QC50q3M77jWvTjaEpiVgBXKNiiIte/kkK3J5iVw/i
yafgU6PSMWwfn6as14iv7h8hHjfY5SMqU2kWy/WThJiiVKrp9H3/2RZcBx3kz4Sv7nR6ETtRu/ZR
+IITcfeoeRFi0M1MCBS8kkLEa4Z8pOGTj6XxVRwn3X86nfonPECALYeTy+1Usg8BlTDKUnfik7yK
4x9Ab6ZYaktZHJIwoC2FdyMYSCoOzQ8uYiO3X0Uppzqgsgcj9baPJsyLizx3H+T8pTz8EuTesFcH
fHoGXr1dXUJQkC8D0uLRJg89+t9668GPEpyyAynp3kn8/BrPutOHsRTdmpJ+07MAEE3Wv3AqiFpF
nxOPoEhRI5M7sBujLVRjY5C28lNYXaG9YNC8/d5ycK+hzdnxuMV73K2abVWAixYPcAkXyNm4w69/
O5yBSdOsqLZh3D7TGkSw6t9sC3IaRksdYod9Ikup0fF7RyNZY/R1xKH9GFGxE2NDQHn5DzbtsM+X
OKan1l7Dgi5hbvA/NZjQ6of89BaJ8Ztr+y07zUibxJdoiOGgznzNxFgfji0+cf7eyhmpPIDRVlaA
93etr05lXzdqTEzAIzeG3Tlo5Vm6wZnY2O6N4MPQNTVvGWermtUsWernQEbHR+mqfRalvcGd7CHs
YPi7BQUcVPT0NOzC8L+JT92vQirFqETbhKgDti6zE65CWsszRq6/yv0KCHQPJNP0YctqpU6XZDnn
lMlNNOYILZgLDOA6ELoKyvYLLKWaRoXAHpIhOEn/Zw5xtCPVC4xpi/HgPBzmD+tYkgEV+mbOpZRQ
F523GTL5ff8LTzgcSIu9FV+scFUFGXazIL3yTZxHk1LUuzJVnkWVEgus3/Tm+88kMP9Xo3pWqfRy
vtVojsMFwxQFiSnndShPAzugMNQ+zFTJTmcW8+W5MwcyXCXF6FDihRgPUU91IJsPMF13qS9mppUu
vCZuHRCFbIUNw93+lVOlQH504LvoOpJz3fJgNu3iUOnoadaah2P0O93USKSocbKxzRDej28/Q9Z/
lTL3Fdqd/2wwIsPO6OxrlLrpaDCWapM01NpGt6Cebz44OU+tqONUf93HCsKyIiY7VUlW6If3g3oh
i1zirN8OwgNxVmTBMCyQoG8iJdCNsYaHpbB/D3VF6acjEfiJSNj6WvXD249feU4wIuluHSueV5p4
i5yL5Uz/hxpHNuq8dnQL64iXUoh69Gbs1Uy/CpEcc0b6WGhCf2iVAAwf8839ugvDLPOHzkWG+apm
CyujZiMD4yJtQysHC9ppbqTfDWwNioxVkQySoyNpJTEl8RBiFtsvO/nCvB26x/CSBd0pPg7sfKfN
oabb+EYdEe3BhGyx11ockzsyfYTZiZTGWIqR2h5ODo/Eki9LnTrHHW1ltfsrSq8p6eQiEDHxnK2I
SMXXKCCXvnkeKQeMFEqr1JKs9g5fRmr2p75He96JwQaHGKm7YhqlNEIrdWG3Xy6flgHSQowBqpZF
KlNs++wD2DIDS+uUjilAoJI3cRJaauWvvsMYC9MNsG6ac9z8Bo+B/YmkojZExEatzCtL0oxgsn2R
0jQQ4fWyqi4GcWgK5xYReFmJ7GYkikfoFt23fSGMOTicYm1rr7+wIrcEPGRJeNf40y+g3IwdHYOn
0M6R0SHcw1D8tQrGETys6XIeNMnoNqaUuXTf56ebitwsduoPnlmiNB8QY8e62pToufquCzi8OKg+
xrUr7Ucybam+0KKub0NWjKS93iQ7eb7lS4X9nzKycYM3vUjkr9J4xvSr9qJxv8tn6f3muGpFVKGh
e+ngjUWC4ZoWgRLxZvlBaPMpbChAmLvrn66B5Gfg6GzxM448o8VvyUcJeICxTwPTpw6kC+cgWjnn
vO6sIUqZX7tSqyGHHqZaDQ6DQpwN1Va/HLFiHwtnTlwIpjtjdHLEe5qU2VWHcs6psOD5TQCOtBT2
/aqTxrc0zm9SClAUFebhSdwzX/FvGBcdqiTCiMuaB0cgZbzbTh99Y3YpseUt6zJoQsOU2a31sy56
kHCjSqSNZ30yY4yPTAW4oYh9EAni6pqzwdP7La/SXsbhfNlWJbVusSVPtglFnNAso0WDo5Sya1+z
6fHfuXiFUOO0x63pqXqYEDNav8nB+WkHWtJFocufANvYKmk76UJf9fBbbDAjoeeqAc3cXdu+QrvG
UFsCpdfMA6B7FL8Mdtr1Lz8PKx+A5uwAz0h7QOxaCnMscdwYKJ2CL6J7ILmtBaXj6BecHyZV7/ka
Pw05rfJDuCLxCDXdbjAs2aLf1SHcsbDJ2kuotnFA8fyZCWgCPAmVhDZ1K7rInNEVlNPvnf3ma3bk
dljmZ6P3pXbxVTQtKb0oLGifKQJgQjK1PX/6jzDQj4/CLO/J0qluVoo0aPzf3AEE3bhgC8XMSPsK
BhEhwuBwRYH96vPo4q9PB0UV+RwChU9rSMWUWVYRIzkD5JRw9SrRXzHiAWuJhMzOQa3NDvny4ogN
D+7M3IbxlCE/EaRf/An+o5ajvHX3QhYDSpz9bppuJLTJ80e0Jqbv2wQHUbOglwM1Kkk3JJsQsFm+
SGMtTneSt/jeHsfy9L3yLTnU5EHAouufcXRb7VNpQpiOReTnAYIJGu4JP59YSesot99xnsVmIkcW
8gNZW1zEhLvoSWylb3cAUd6FSQUDlxLxyQw7uBUt7VCaI6huQ3pcokKuOccJ+raCx/xlKEw+HrNX
a08hVRRXVqCnvU3YvQ6WLjJeYKLuMRrFPaZjxIRuoY1G4okHSU+K9br2Z9YijFNqpLFTF8IBMCfH
+VTEnWJuK1e//WFatZSkUN8qeRO4mWqGBoQW/0DGnVOGxSZNctsRMmC8DPzLtNj6UY+GGkrOyFc1
hT/4z8IZ+LAfyOX6qkckPAEj8Pno1AtEqBUdoeVcG0jeQFFnncBv5hPHvsciLHBJTTyrDCPADJXH
Qkt9fzd0gt8KOIdIrHb1OhBtsU5upCbWLgMRAHgLoyeH3ZYPHYMAQxoctm4jxrpSiibMPDUrdMlj
tPUsvFxWfNYYYpdx0cas8d4Z+3w4UkU/gItHboVV+MDUgUdDMggDFyMLx6sF7hW4sN0RKbSdRTPz
I/kggnQ223WwYOSvkydt1joZ3XUs47sh1LJtcPoo49v0TT0SyVzE4NGACXhtuHgHJWT5AVjdU7oF
mcit6zzM6QjFpux7/TzTrmgx8B8HXc/Nln5/JEuwwoKj6hhaZruh04FgNchuHsx45ILB/Y9blLdx
gNzPpJQ+W4MjsaVuNd2LgSFlvLTW79+MTdrfTXTyYg/sDL5m9rN3L/yj5XcGEnNpK5mbrEfP3aqL
QgiTKqBKMgyKFEzbxzhZWU0ylMwnDhdXB9FEqk8nhyZpaH+4Y9SLDRmn8OVY4+UsGsNEbcz00mc6
wfsQmX7Ku2KYOwezjCtuwPnG1p2IYfq+CevHsS1OrUs5aqj9XX3ickqPXENUQEca/oYDCjZ5w8bf
/AzVmLIuJqaPeL8h/jh+CkXHIPlUXlldCiLETBXWUcpirQVsBJcSBMSqlS9fK0PLM7RvzlXuLTuU
tE11g/K2qVkQB6zz5/V+X5CFrCGReMzE2j0ZS+rTOPpXrIcMIw/ofpke+U5ez7xfkhdKAO+nff95
QySsTSWbU/D66sGPpfF9OH0P0SEaKnYGlddPFuhaOAzaq077BbPhmDLakGJbyYEGtPWvXCg1gZvW
OnucxFkvztsJjZmZStG8xhroCFjyDl0vZzkhdw3NGhc8Ctc4ejVn0l98s2p3qmKOjQ7w6ROBe9i0
+3QPnGKt7KqhHs29zJNsgmf1Ni2UrhRFSELzB3IVIMORaFTDkFp9lSrINHXINShRFZVbKmT5Yxgg
R9b7M3CYOkpcbmtvgJTT6BmHJDy7PzGU+34XZoDqs3/Jyft2A3mSF4V775K7WY7gwkQq6IN+Xvxe
nHhTeWXDjt8WBA1dCJwJQtEs4oWdBD7dUk6oPp8Ag2WmDHd3K6jCa3vthpdKMmUOZyzZfL8tVDuw
4f1ouU7NyTHHUvx941oUPIXYRWVu4F4OhWv08LOC8M3NOqgNDUSZ2qTxjPxaUV7z8fffjB1CgFC2
6PqF/a3Ieb8FrpWvL04X91IUhIS9CmWOjwXjl+zzqRA/kyUamsHRB9d6WU4aq9xdb+oQcICCSFbr
eC1SjH7m6mEdzxCsfoMSXuWanxzsis9bHQXsO+LRpGZC83bR2ONqZ8+wpAdzKjchVRTBkE/3NoxF
jy3/jPBy6Dato2KCB0S/UKpmsrBtAiEqD+cuM3fzq6yjHSnwEBNPSlXVwFCoduqg5DD6DFBdO1+y
JJy6zkCfwneVNH7r+2/G3VSRwSNdvzFBtLR5CD1RJ0pm0eYNp5H1AdswPx8wriAZZWH3nyc/xCQ/
4nyX1QSI9QXPBCAZRMIJ5P7JjX7ok2snFA7Mw7NWBKxti4Q2Uje3ZTnTZM/QaczXFvMsDoht8SkL
hqiIACgcl1I1EqCi1UlouP4FN7MUm0iIQsKqoeTDbAlnIGzFQ2uSvNp8M6FNXXrr/UmmAXhjUT0t
/LahLJbaM2qBifQ5ZWi0u3yQrAiwrhL9mRoduRelZv0GfrsZM5IYAdQKksHzCuVvXJuPkePM3x3m
Ij8KiX15njEwzEp0x0FLiIK7Jz7LhaxIcS0p1D5n+lIjbP2qgklCn0XUe8h/xkmMXMRWjE+9Xim1
wfmknNij7hzBsaB3RMwI1FMLsbI3Drptv9WEOC0bFxBnbjpbI+8fo6Fy9/TBR4QhELJE5n8I3/2e
2R9dUp+YjWi7Jv+CXBSgbMFYD2Qkx9/5uVYQhhkDBrnZCeJ8rnR66r8wihHt9ES5fJMy8btBzUdV
1lyRTu5CSrHQ1yeB24tuj1VLhQ9E1cWX1h00cM+3FvAEhrfl5JaW7STLfCm0/T6BSAzwnFm/SCfm
1k2rsvPWuexjfEi7NylFhzME03oZMSqKtUInVslWAVQfOdZP0DSEG06+115csWU7mnfJvW18dpKy
8sSyzbYs4b0DzMXi9ipy2+XYcTeT5xCo64iso/+qUFpKt4b70B9u82LVuG7k4rrmg7iccUzUHuLl
0gChCAcviE1yypidC52EVo6FE8A7OU524gMorOS0KN9CG0aBFA85dPMQnS2x8FxY0UcXrHCQ8NfZ
QiLV72wJQPNrhOX96FXzIbjQMIE6YdF/MZ/qlXK1DArUicPPg/+/9Ih2yLzprGKuMoCSvihic+qu
JaHdBQUTc/6KMLzPpdFQ178k8y0WlTQ8M9ZVU1XXU42UlGzmFdwiC7PCU/Pwv6J+hRulQVoxXDSp
iKpPzW5k3snnhEL0lc3bLrB9gGrYBR3bVkINY0Q2Q34wl9qw6hQEa6bxBaFbskxL/vCLQ7S/wdHK
s1GFLj9mr3GM+MftDqnTH7mfwXtMmgZnSrSrKad5E9zKcwG26/G7GtTZ2zBOWicUSQYfbsTFt5Iw
D+xfLTlI4PZSmDK9ef/YGIuRLaO5kpYumAsEKkcRjR3heYJGiFrTKc/YMx5Pc6lD4YDGg1h5ZV7u
deQ/sPoC4IvSAYpklRKwMZFY5U6YlpgROiqpBrBIHQewFAAcf+KI3KarUTlg1aXcw1E6Sq9NFFQY
EVtfvsSJihW7mEVkcXqL7Rq4xBBzFyQRpuZhTvVGYm0w2uf9flgizDLh7W5adSaFjFYHKzwJ65Kr
fM++pHw8FQSNmLpkT6dnpTD2XL5+7g8jyQV6h0GlEMpjqSaIO3oTDL7Oto2ykzFdCwEMz6sWBb1z
NzVMBkgXtBdmmq3vBmxLtbYtySHP3QyRnpG5AQ4SKuc9f1CPS3pw4pA/7yVKYsgzEH2y7yDt1riz
hRsl+1q7XACFqaLRdBj8FATX9ryVDoAgmTGgw+acqJkAj0Xgd/SugD3zn5Zmlu8E08GkwVL2EIne
N4cyy/0eMopSn02KpMwIMaumMMtINa85SSVOLfECWFADeSa8mimXGJZe3FkVHTiLyfe4s0QnJ7WM
vOCcY9KuxoC3415v6NFtthMha1TnzPc4TjLMQIVM53nKSTjl/NIKbpMuzHqrNWlhV0ge3mHI8VHB
YtxUdrtLXcoquuGSsmco75iAN9bu7UYCK2Gv2Xdah4zv3ZAsQ7YXtN99rI9Qz40yN1g9q7F/gHn0
pNtYJyb5+ZS0eXiY6Lhxh9IIvJW51+YRTWsYJZYnnGgmDTWmB2+h/CQoFAhAZM89id01HW9oeXGl
tzbO7tVOvRkWECv9SLLGSSWuQAizHPHgZv7DLFOVe9WPh50XGI4gaS5kgQHFh/SBRQWy6uRlPWEW
DcQ7EXa5Q/q6G8aFF/IDVODSdlVSNMcXMDU5Lt1hrZF8x0AyyfIEv+IpHRxcCGkgVZq/8V7MboO2
7if3V4tROdKs2d2/vgbGYRSIHbpcQWp8bVdNXfmhGR/n3zwj5A1KVB2lAt7x6pjcgNIJWxC54Jvn
z/wiz2WlyHxkYHg5D6u0oaGrfoMZECs1JTu/GzjqDBN2osMGYecSJR8pPZynS3wG+E3dKB7lwGyq
28EUxlfhSTcXCPcuPpGq4Tj8Gt+Hb1aGr9uTAaMdKPhfwCZNQtR4Y3AFsdBTFBokDkoTpQ5TiyAi
ZBfsLlZcWVcve5O67mMBLm948EW3FFcxHMuQnIyvt+2jBtpBr8RdJ6cuCEh6bBmvWE8xovWxAigN
nC07aZ2V+ksTntKeqOjNKTOPDhAXHRk8XlYXRzXurL34aB4NGpem6xruxZFjpS6i4A6JZglgKgEN
pBOBV6qUrBvaK3Sa5F06yKvadLtNdqwK+wK5yOHSOja30zT2iD5o+HdQU1QACa04AB4wKsQyi4Mn
kkDFWxezwtYi3ns2e7dqtSR3degebCdLk39FXXVUf1PlPwQ/SG+6k1ah0JgD13BE7wuvd+S2K2Gi
ItA95qxWSaSz6sv1TRmnWVcoxEiJyxA/4ZYRRLV/Nucel7mAcS/AFYTLGUnpOFNXMA+MH7bRJRv4
kpzSsJLRlYk6cLQQJW0fe+MJ39JLARcx3KD4C1xEX8pWyDVI642/egzolUgJSjZ3VGbGe2Rf4ndN
zVA2CIRgHVh/TgGge6RPU7mjVFB43oHUQylfmkyIo5Hbr/KYjFq9OqLyC9RRYHOGv3Er8MtFiqiz
LBSvUSCyaf9UbbN2oYy7v8MwYSyA1ftcj5ddrLTQFPGBopN5A1fxC8fJ7bVgnlLCwiodIlyNd6xh
kAoDMlNsel/Y9pzp/pyP7mJIw6htrKQQWC06nPbeJCfIdFcOYaoVmQ9RHB9icmLqhrntK0n4Ulj1
m6COLB7iYi0jZf2Q5+/xXSzMkbFmJ2alubXLhAmIjsmeyMmyvQuFBgFu8B+Y/aNGX8VNnOLrCuEX
FbXZ9wKz9lywpotZTnCcOV64mKxqY0AMNIQHWIzVYLJQA+sjILKw9hiW/g9NYOcsxMEY6cjsAn7e
NAnPJuK9N47XI2VBRqxdEMyx3lLWqTNjiMML/w9Sv/lHevUrzi02g7ugUFyDMVfDoKjEEVaVNv1g
CYBnQjyJgKu1CXjRJ1vYvEMVv8BXPWCNlCyndfrw4YLcV9XPduDWauwYmjgk/yb+h2+ev3h9n1/Q
Zr3KvWFFvMbBV36Yl9YC9gBIGDjdP2EfpFdi3TtxRE1zRBdLThtTEG4iK8nfC5eLHuFuGwhMkXQR
sllv+kJVVHG4PR9/kQX7mknI6mCqr9vsuybCJZeUEmWFZEQ+IM83HhtU95gCVI83Lislqj2k8s7r
5yRL3RMquE19q7kd9B7eXSTMb09GxyMkJTZ8Us002DjOrv8Y05Uqy7g9Jfmg4YScklztVJSaWnLJ
qcQxcjj1FDreCoDl3cur/3y3c/k7zc4n/73Hy1ZVqZQM6nI8TgwmgZeXrOnkl4TUCfNpe+yZtGhk
CTADlxx+kcIo5I+PfNbTgZRIuAjyw7Cc/xAKKyaV3BI3HIt2owSnvK9lGohMekR0USqhmBtdNkGE
TaADhXsCDsvAJGyHz7ZZ4ghZEHTmUK20MiP2rWje6hDYa8gjs6Fp0dZyhFk3NVeO2ZzreLY/BSyU
Qss16VLwVPONXFGyGvrjfK98KThAPOTgE8ukQYYlaiLponZmde0sc8EtvDnBd+EvmZte/OMLIAN1
p5KhyqEHjLlvb/uxZeHkOJfIFoRuOCv6LnqeY7hVxA8QBXTuKLGg5E7cJUXsUuxCoXYqpfC/hI9v
oOx8n/3na3c3k85yIWXXdeib11i3/cSob65zYEu0/BS0ZTGu/zuhop0yHr0U5CD13N/dNvWWyWGd
NBDQ8ISv9VvxzuHzpRvQJH8xWNmG0+AQz07H/zTiOSlJqTZD3stQY+cElyHoLEfrZ7og/43TtGQA
1nNnWt5M3hev36Ojbu2QTUiOeBwOJJ6xhwjX87UEESWuiswWSR5gkgLmylGyHHNeW0UIU3Fw49u8
T7/Wqu2tTb/unyZo2LcVHCbofmQmQPd3b9AIQ41F2TPwuxqbxS50z0tumdo1GWStQVM5hVzjjD2K
tzhAjYcYG1oITCwUkaJLxqaoN7NIAJ+QqBuE/POzsYk90HKvgLAx0fjbKb2JB1kRR+kPOOpkspCf
TdP4YMjmeIxEXHZRYllfor1+IeX3L+F32v7Kxj+wWu+eaPlAF8BeyZ8JXfRs/0TMwD5281zn0Hwi
HgPr7AMdvZiqFdHZRaeUTJnwYw7Sv+eekLKeepmn0gro5FylmMJicpHuRKKnFPyMB7Seaxf+mQ/I
SaGsIePCOQSLZ3Wf20p4QDNt0vj9Y6gDj/X0iD1OLFQKU2hQRnf06pUMKgBlw25Dtq+xCfxUksH5
9PBFfWev4TZSAC7t4Y8VeUAKMZyHYzuvSEr4fEZUJR93m1qX+bhaGxd7oPfnAz9eRTWynrQZ2ZNp
RCrv8Tx8qt3J/u7r+046ZSXReUw3ZLLgIpBeXZVwzFdU4YTDGGsEGd+/YDm+pUN+mwNSAFy3plGt
SDwSVxy2M+OU3mwPU23EHnPslPdliajUbfM0D3xmvyLp9UrfKC3l+aNeO35P4z8TMDDfqn8OJGlf
C42TSOM0NO65ok8PAKPVKeyOW5sf5/o+ZWLx6ilvgm+/SbcaLuHIqe0/Z/Jf4T8asaauK2oqYGUn
X3QOYzRxGA77cRug58URDo7XF79KPEMjCAQaCb9LUb1fvKHxohH/tVXpR0yt+9KIGCpKdXzJWY0S
qm+nvO3j2pxaIGTgRzpeXEvisxKrHxAJuKswdNEGzJrldtTVCC7Kmm62wQjoOUbXBzQPTcMN+ujG
EJCxpO/Q66MweiyRsIarfWK+2YhleF7QQsLfaJunZSmBxCmzuC9/vlmFjZup9me1CT4BGvpCfhDN
Hqxbb8hw4HWKih7gfOzNgs3Q4/7fZIgpDxClzAC/QDM8lEJKP3eXRdeLaGiIp2xcFS+noGdNOkXY
90NRtUHmrYAuzDqDtLYHzK4pXXCO7lBkKG512deijpnoeACnAqlcD/RbYuiltnJtcJZToLZC+mOO
Dx5duZJSJxuTQwKVU2CVNRK2H7JveS5jL1FsxWFWyht5UBlMmgSN7ClJ0FKhZbTl9DSaLUa7pq9x
vzbL5uc5/BhZ7hFTSbGaoNsTjVhHAC55kkEI6dxUYEAAd6bEE4HWeFrdO5/vdGpahSLMCrW95wj1
0JozFG57JXikmi4jRYBMtmQA//SXZhFiofcndTHcohJpBclQj1PzbwKVqfHl9k3Z6/vH42JLesrT
5QAFQoPVJRkV5LusegyZvygRg2zMpFWAstpAqkntceNiY2hT9IP1c9QXTTkTrr8eawV7y1pcbr0Q
vdRTLwctpzMHexlMgGPNfrWkiW1pI7muy7ASp1YqxqtTsK21A3Aq6fhbOqByC5RqybrwOmuW2sIB
NbcHYZABitUBie4LYuu0d3MX9WfjenmcLQKeEf9srq8VGMCx/rUdlYnDrKCcl+HeeC4obB3bOw02
yCTfLwTaDkZTdnt70esR2hvZIb8nFhePM2Eh5kkWB8wu8Fb9lib8zGhKJxrRpwq19oZqnrafz+ze
L0mQhVNqR+cT+VFTcUgP+U1fHGzebDzRqssn0YEZOTun7hyL3mcw4fkMWAnLGYXjIJk4dox84+iI
4pmEBVutm++cIro8/TiZDOl9czVVujH79GEVmzbLlndlvMU+yTDVGHqOpcp1qabcxgT5kvRBbT76
0UkMn9M1WyBDSMRH8cZfV0fjeRehzQzHS7ZYueRKQ/P0eFdL1FiniOsKXU7/ArB58tsaRMF/Jexb
vbWsgq35EndeVDFQ4BatJ2rEbS/+FTXQiX7cAo9W9ELT22Sel0uZCPCLZfT4h/Xqt6oxaoeIVIt4
EJVa1dh0yY9vQGtocAySyT+Lx1DLbPCQDxoRTgFB05mYGXTn6VWXAy9oNVxzgvFqUcpX7yPCFgHX
LQ/W+2ntAPLQmwosjfRmKcITF3IodXqbre9hU/pptFI8LWOzeGWgCWwfSmJaUcX31FWFnRMToRgr
tOLglwSWyG7u1nJg/ZcfLsiqlczjCz018L4XXT1WmgJw+NdDhuDE1axPtkUYzJ8sAf+wgidzoMl1
N37dj0vl5+M1Q8Z1xee/GayYV/gL4nS+pVKGLXNTIroZMwMJ2lbFEI2LmgNSQpKoWvPnyKzQHum+
PqizNs5IOvqM7ggfk5kCl2Sr5xiTg+OfF+gS5MrNTmdMUspjXhgKF6kWqMFFgqQuVMiEcvGA0sxT
mybS0C8zSVM2uTpdpaJpo4fpGSyjCsY0g8+OjLDAvSuFIiOWPD3QrL6CU96t30wspjDC6Q7JiviF
0Gq/hgkJLPnMjJm4JwDTZSrp1YC7Y4PNYqswN5IIP21h7gHIptniVhjJ2EXPgiMEIkzJswtM4i3k
XLIfF+5DF/kwN9wVfH/ORhyUjacSLjCJWU2nafoQPYdBlE+QoBnhZb8Su7HqJr7GyviqV9T1n7uE
ZLPZm2npGFt5VJVj2XzvDMEg5tPmbj7X80RR/Bs1AbJV7M6ZGQq4jPC49OkAZY8xYgmwxn9KFoVb
Xk1MTPzvC9tPdH1JeJAdr7j8/omfFY4ONsglKiLJdJisjII/yryX/C4NEKQNUOGImOHadP86Y8xf
WUuwlcN0Iyyo0ZYQ3D4+HCms+YDS9Wz77RFia8Jh2HMc7gcSkW2UzmSRlGz8GvG/j7ca9jsOiHof
9xn5W38JdJwB8haw1DcZE6IFJMqB6NygqxUGkjmi4HDo0AdAUkDiDykQEbOe7Lou+LEXoZCyx0hC
6/6LNak2mZ5fSeYATJKCW+jUIZFfCNGeavKGRkNFhM115AlCltHa620WQcXekKz2s0r8YyuNn3kx
7Hrrr8lYUBKDxE17DUMF79VEIWUlkBamtsjZFvWf5izSN7lQgeWMeA9sEctozQUaQUEF//TECq6n
5PpJgIVxp3CMOKAHRfUuePBTRNZjiIDcic0K+2KQJIvbwq5KuGUwJnmuL1ob2ZbAZ31yFjILba3w
zZknYBEETbXQKrzicNyNTWa2sE7fsLn3y1oZO8/yoX9gBTrPcPFA2qfLvi5M21V15O/mvQsbB3hb
9cXoQrQ57y+JxLJI2Ex+9iFZvho7N8iItVVZXGugZfJNjLWz7vlDD4gvxabA+qkHyT2kqSbHIp8w
LnB+SBsoyLWqrKPjIup6xJu+4dUEWTAwAotYvNoAqA87ZogGNlMlBY3dGoOXqRC8D2/lDVwb+4X0
HuWprAlZeq80yatvG9pmgxPWDSVnCkrdPg+vP+93WqqdsNX0QRM+DBPMweCY2CwpGIwVYvS5QYaY
BMyYjkg2gqmWOl+W79bqIrEEz+Jbywt9PNdyEVr6oOZWiscjQUGm7aVQv274aUA2ucboTw/U1a9b
YtnfmD8OvfIX+yoGBZ0Z90z3+GipxrdLX3FO2xWzn2+90tfbha4AkEYIV4JlYZpwx5mU0beP64TO
sRRr9chtnLVo+EzEi26MwFY0DmzietuW3m3IC4wBO4D9BYEWw90VAsp+bHqlYofCczYlDBoGfZRw
g5b9qW58IgDkcS6GYdVL9Y1vToddFru3jLflJtkULNZGg1BG+Kv5UrqeSJPCFOYulDSAJUk+Xjey
FqPo5MyI0wjo0Bh2ev4yOE1YECFtVYZUbUdUYxizcdiZyPUmWIt/DcV/j8vLWahI/KwJt08OX88h
TA97i4bQ3AQyYt5HGWNCj/6XKOVHqcR18jotfamSdTi6lTGldYKNJsONkBI7lrR2Zbvx4LdDbxXE
7sctp5DTZnUoQi0X5+E+wpVBcow6Y19q2UDoQicfVJOVZeAhxKvGArARqFYy0qO4sTj3roHyCmUE
RjOQMi4535jJmiCva3QamZcoVhGL+oW7WLx2b8T6mWdy5gkJFLqW9SPV6b2EOQcAauTMn+8UuqA/
bL/C9j8aR3XC97UZ3Z/fn6oZSVLWJXXCpAujuPoSor8rFHZer3On6i3vs2PvBZv026+l/jooXKn4
EnxnU0ILvZmNtGsn0ubsKLyjGkQXfdILSH0KenhOFjYIfGrz4vkWJanbfv54fqKpVPu9KALWSlrU
Ul9Fdon5YYq+dr3Mf+GkGGA8wchy63tXrm80lhcfsxDXrr3hm32BR7yFl20GsNP7lPDoxWRrYyVX
PhOBJDCof3SWRxAIb6yTQzChktAltPZ5yAwDlN2TkNBmvLiCMh0Iq4PzTmY5MAJ5bK8u/2DtTb+w
1K+woMZuL+9lnX4mrXFe35ml8DXYvUg3TQQOfAOQXc4M0FzUXmnd7P+sd/g+q9TEqIUl4+4bibk0
TllqS42/WqqWq5tFgD/J56ZzjByUKFFdw3X/wPQCAZTusiKZGBE7KbyYEbzmgtzSRyTdtEipQ+KP
YXd5FiUF1NkN8CC+wg9safXebFl28/HVBEq5ZJHMMOaz+qHzqccBw5YXqqa1K4c3nvLDTyrhoekn
4dumZRH+1mBO/jH3FFQ+tsDgX22tSNpiNjcypT9i+yMY4a6RealiM/hAoJRcDO/cNBogJ+tp8WWp
HdpzBF1+RWM7LtSn/kseQkF8hZewiE8dN7x4I3oJ3f4HUGD7lPLwDOgJb2YFFBwjxJEMCGxOgj+I
Zu8adTND1okeY39tOcM2UpkdQEv0CrXAv8dS7DyQy1pgBNuESZ5wE/cOrN4xzgdn+ogkII9wQ0z8
NrC6CDdzP9OD2xgwJrXAbnzgFyT2FS4+DuFY46F0CTx19UsSVH6W3P5jD2svQbKR0WSZog3YOeag
HVtVFu31qrn3k4x42w8pdldziYVa9Mmj8QXvmrBkiRxNhJReZ2dLtCD1fbwQuNMzEs49qZFboT9s
TtayjHhKia7u7QtqpYzxxNtzEoFWNcXdtUGibYn3KNjgyWPjNuH/5ffmUkGCKckRgyztuZfDC3aV
7jRkM8NCAGm465opWsaU0+ciE4BUFCsCR8w1wsWRm1rTVpyfRT6SCU+0y4yKDfOONn+odj/+Pazn
UQWF0IUYSZg3+eAnE4jBTz7fvXq291bIEoDi4aix7LcS2D5D9SpErX2tHuJnHEFvf/Ii21rHY3RB
YqNuBpOiHUWuN6CLuVqMprtvuJNd9cgJNPg8eedGAe8DWIZR6BdIZPGTKVoIezyJdwsmxW2xUelk
AgGT/3zF/NUgBzkansAwBA/ytfH4/743PVfj07x7xCafI3IFImxz7Zn10Y+uu5n3diWuMo+9lhkS
PzIqaEyPJgLkIpMyVYGKb3rsO/aV5p1ML+4wZlhoBHNu9ZMft7oEw4EYuKvTRvhFHpSYAf0QXXTS
9AOBOaNBMnkhtBVl5uiufRXn+YMCtFEvrli5x1SIi1QkoZUPtEAEsOk1NIYJXm7Vb7S4qAhd1Sbd
6nuOjsaf3a1RL+t17LXgX7HdY5x6s5aZK5czN4E01PII3oMVJYOROOa9x7Srs2+3ckiKbRMPIrq/
GMEORa1guWN6fbVnw4LW3LQect5yrhpD946N5WrtxiobO/OHT1QITDEt140hKsupTUvkXMHehMGY
iAScDAbUsSXM3PiOubyOhnhfeD+zSvcKxrNcp7OqHnHBOsR2D3QIwY49Sv0BWMxuvkD/KtHOg6rF
n62QLoRYMHKw1U3DXEM8ZbLybbo/3rsS++OyJeRec2RLhQ5e55VVwF5AWrKDU9OMHIlSbrJP4Qsi
yNni0IlQ/UcXGGyl9+Rdj4CcGsn9KoPlGTvqiWMG9SJQQ6CNBMWK0lt8UoKoiNfvy3cj7qpSFULA
C0XVqJ23B7etH7qSg7idoKZcZjj9o1TuiBVridB3Jb51DdpARdDh9QTcx1fl569rmFPu6uZdqWnC
+OTbeultViaXZ0tXKDGbPR7hDqEgY4Zz9LWkdMQqRldPJ1JebQ5JNdtSOeBTPd4qt0vnty97cR+4
LGxGQ6Zui+VgZ4rAiCwsetu/e94H0kqlW9U2KDbZMrHdddfIXz4a2fQ8nOvdbrofe7D36PzEdErA
2a02LTqeVcqmd7eD9wdL89IEkTZIuDXOAWfhWf92aAUMEhJURG5pkUx8rGHRDs1A1i6h5Y5ceUp+
AqLZcrMCyK3Yea6sTn+rWVvnMBuTUWU9jf6AofDYvyCw6KtcTsOqtoQ5h3keEIKbAT/jtBjyleZe
ESTFW0v9JN79LXhuuxwZnnWPC6PQRHMqIyziD3/O/dQhHwmUrDZSy+i0IcuY5H/8sGvngcGbs3Ef
W5AXMQXuYYt/3VhlMh0PAhecqqtgNEHSuOdk2EMK/a8TGWGV8eSoMjqxgRsoNUUaVUAYsq+POWLv
B9jZJWXoTrX8jnrm0Ex+qbEIJPAofdzAPC4lSYHvFyaclOsHlSXCu10jdCTfPvHoqoQqD/aYHldG
IQhP1qtXhvs9s9nMkwZf0dhDyIsFIueb4q2IlL1lH5MM8buaooew2dP7IPlJaxr567tozTHFS3vV
QR3JAcmexGtdO2MW4NZOHMuETSHdUd1k+OPr6UZ8p9zjmVIHy2y6NsUpN5aJLUfhZT1Qdp8k+giz
E4RZku24GaAFG6rvi7KvutjSYb68dtwRApAFx+MhB2Hbhk8f9QgUyXAbhVWehCHVNs9Bm3hMrolk
pjvTSg0SlZobrDmmakVx33l9NJJS6BhRWX6/DasjiiXHjUepwzhdSWLA3b8CSHcV5R0jCxKyHILe
vTcVK3KGDOdoU/gnI3d5WDFoVli+1CV9A0pyDzOGCnKDDNr68ZMYCtj4HCiJ7RHaJe/AxUtffmf3
YGfXFYKzTMj5U0Wh3Ne/+EK5hoCqWFCFw5V+ywYNw8F7R0RjvEl36YNwIgFRqgWpm4KDQlKmv3Uc
lspYTtrlo7wfSxtlYIuQZYoQYWZKDnn5FPTLJryUnAMkqMRTE2M9DJYGHpu+J32DNhWhR20h7m3d
k2k1SjSWrJjBpNurcJhuJux2zoPa3oJnOcsKlaaVyDoLJyJ882YTkpzisMd27hBdB+9/zbetyEFp
NPmnhdddo4bnZjXp8oH+qcXnxysW/LpqAMt8i0VeSsqc1FF2BzbCJAvrS6urhFKj1p+EgiFQ+PjK
fOnsDxOphi0ku/E0i/ifL4jfdVfrzT7xd30fmYFLW5GXNtrOb+qYU79ydwAuISRELYPZUVzpZZQo
PnXl8aaiOhHFKacvFUT8MRxeB3AarSOdhsJC92ARDaoPYginJbp/ZqoQbK94yw6EfhymDKdNza04
kJGhp4SbL1+Si7fAa9h8Vc/GRBTDtjUXN3h93U8k0FfUxkRd7U+3LZEKU8Jr39IPQLvgSJuVe9tz
2tMy9V6L3VjQAct/lfdaCHCe0Rqz1GPrL4VbIOuPjhtXNDAB7VaHT3UhUwsGlgZ+t0on0Cff/JQq
T8VPB4BwZsGzfH+w4/nQ6oLoSXpesboi8QzbWc+7UNn5P4X+TUA3vPX9IpoCcaCcn8AtJy5sXt4t
zey83uWKUA7dlHyMnMhhQzCkXCFVmA9ktpUvRRdbssx3g9qkEKj0y3KFfM4LOFy0ZkhmgJIdha6a
lBqBjU5jHgofKQu1BQ6cONb1LV/zO0ktW9asnH5U3d76Eto8hrekoCF6zx6qPA4OlxH7ws6xrd1S
zPGQLmpn3b3nfijPGoygcQpu1Szj/b1rEylp2wOVqXL3XKPSuqFLlwJIcNTXxyHXGxJU3yY6xM9J
p0mBgDGjpN397hKb/RIhXF0283JwGUw9HxsPfJooxrLPYqEl7X+fTeh0dMcOJoKPolBl12WHacpV
hfLvNTu6ujXCl1+Ss8J+WbVuCGlnITCREW97HSFT7o9d4YC6E7rV7S3N3j5TyzFj7ODjVcHMTDTL
RiV9ODL3tZc2lZM+D2HOlAx5RHOWHB1zQMD6VkDweSEt6lZu6qCuikAknpNN7QTC6YXyOP7IusJz
dNpB6Sk1akYQ32Z+GOvGUSMoOfK1A72Mg11qnU+ddyPTahVaj6D20Ai6XO0kVK4iBlLUGlbQhP+z
pidN3djQi7g4LFFrTcHW5SgFlf1fHyXAlhd0I6SVNVQiXtiKAAUmeiBZ9qh/Y01gx8VBeqZvuZ7u
bKrMaigkcGfXzbGKcd2n+xNcJHVN5lBNod2Ai6FdMiC1YgIQI3XbO52FglzjicdKBa79YaYVUJJ/
nspEJru8nghDuzVSQ3nL7kW/5eqRevaf3gjQ2IeSiUc/OFaAMkl2STuLA6xpb8fOD0kJXpX8BC5N
GhSChxKfbOAlcWQmxem5dBi0vpwv+GSJAZJX636RKex7REFF0H6SbVNBdJY3SOMT23AklzOssZLy
DfllXnYrh4p2P50zK960zGAZlAKWQHgFRxFcZ2np+782U8sUO3LYbOq+fnMOUudBNddNzUFi3JWO
Nr65s6eeZsEtqc6SKUebURSbcG7BOBIpEL64/f9bmgOZXhbqve+yAn7OEnqKWv33Vf8GRTOzKFqS
Z4JxVmbqWA5REYqLKPPkhtWFHwQEEmdCAGAK+WPgSYezRDvR6VyU+Ksyx2VaGsFVzvIIVt+D9Xwp
TNn8vd1bEz62xL/2MdrxmJVhcIO2bvLasP2zMYg/F2qMaMjeJqEd7h/sJ2k77yCKUrtzaXt3wRLQ
y5HtAMl/r+7lnfn2p8xFBTL3Uk4MrLMZAKGRFXZq774k2Vn7psHNao9L29kn4JvD8E5YiUgXTaAd
6zraEfllw8k2lURRXZo/NUT2EXFhkvNxQZeucppk3Hie2T3sOere9DO6Dxuxk0+iZ5MGQcBYdstJ
fkdWD64TFd+DYRz9/nVqcIJ1BBFx7KMT424EP3KOF2MpFlUNLe9y5H8rBne5/yq50Mo4mG9dNNWK
KCAL0ZoR4+jpJTQ/xfLDBRfnKZBznfcmemTJl7+idRiTP3FoGz1sivcQ1Y0OuPnGRxwX7VhSlk+2
0ef6w75Vwy4Cja3TYtpOHZwjcua+FEEWzmU4G0hvwwAer0sTSc1mXejKjA0cdH2ZoIoRkqc394FS
shJD7oka2bOcN47GCZM9X6t0QDSmCvsh7vjPKSk4vnguRwI4d3cu4AlHfI7ZyR8agRW1pmbC4lci
wiGrgPZPtgYvXXiMD4LDLIbXQpEe5R7YYE150iy5KmsRBAp3waDx5r789z3tHqLlg/4YJah3lv0f
oMfXZtzAxwchFye16VCkat9lQkiiYaF0aDscAhm8v0k1N8X0HDQlEWDpwb2yh5RCumpAXLxcqpQM
/x6Wdb8Ku9IYoaqZtUgFIEI8A/hF/r13X1loU23MZMYD66iGm1gNBEzcHdFHasxzYixdkvJI1Zqp
wxwU+mx6kI0v4p54e/wyFvKBUKhJY/lRybNV9scBLDX57NH8T4Q3Gbdz7oreyt1f5lpi1L5TuvNF
mAiHF846fqsqEuaUi2vtdrFTW0t9Sd1Tkaeoakso61K3lYrN3BbBu3ADtGzHPoRVgnoQKqxYZvzd
KMwHQe/fzpXsWLGuUlfYMiyNYaPsIsWL18bwiOkNxEdAhF9QFKTKRLtpMXFK0/CMIV8S/Tj1idra
mFSQolaicP5KwMDKtR8tSjKx3BtFxJ+6v1w8y6Cjine4cUWg/n+/QhlltVJu6j2HBSqQN40yKjTt
SbmeWjoXHlQVPgoWKf1T0xTdj4/AmozFfid0b0alEVPMG1mNfUyOeSVpfk3itBV4mr8Lfs1wC2sM
ntvXMScDRzmED+Yoh66554051uZhDjInEbX2Vu7Zzy9mspwE7LznkOwqbMzZ+SmQiIN9FovqDGed
lNDZwiQ1L4V3fS+M5DboB1keLmwaexYdTLrvMCOm0gO8aVAe32oCVyUU8VvrHZc4e+H8fP2ghZB9
cSwB09xsK4xrbvfeLFCbJOMma+5D80ToCIjuWvHahrrJjqjHBLK0z1a9MkgqqsZhW3FDECBlppmQ
u7RqkIFiLnZr9EgVnzgcpoBVBGYAQ0FJ1kwTLjvG7HwSfhqHK2eI/NK0D+Vy4lICQV4pbO7pFgDJ
z11tws2aOQDoSzxIv8VQbwFRTopQS09ycCBkDu27H0k4Nr3ySWT4teIV5Q5Ir2Wr1B1TKsDrzcLJ
xgUn82bsNf2UvMRXYx0RImWuTSSH/Eb4CbLMaGnkr9cEQ1YkWz/9lgASR5oXm+ESyFpkH8Yc149D
5c54wWnz5M0yV5f9o0olqLXJ7PiWYd1oqq0tgdUwNw94hVJxxDJfBlAPsrPywHR9ZoB0JPVnaqdr
3CgR/RxifGSqq/Zm+BRdGANoOOP1F9kK0sv0/0/fHYv7w3SzaE+UvbrO4SgG1VBa6uKSGrqeLyAu
ADukjzeX6cYycms6/oPNF3tb+K4BHc0B13JuA1RlLlXkN3wjZksUPVOYkGGLsbeJ+bYQIixVdpMd
FnIwCyIYE940Sj5xf+drTkEEpoos8HQQInRSK85hGTgMxbUxX0BgSKdm7v2PqRrQgWLnaLRb8Oo7
4usFI7SpSckuasP7KafzNLC3rS8GKf7gvzcp5iFdzw2Hm1ZmaVvByzGUsato80gRiGsapczmsolN
EfcPqMa+SrvfopORwcewbuKGNQ8ihyThHuWxxrCS/L6N1P9xCzWluX9oTU2RJciBoHEWBRUmdWmG
LuY1Pg08g/mtgFC+b1PesvLroi2UubmXUxW46sSLg3+AVE2AALIs5MkZxXV+B9MQBU8RuoAivOir
J3PgzhVNN9teYxDiZFIpJUpkWZqeYdHLMeL+2qjZNUgzLSlD8w23ewDoCRu8JZrpfUQ+LmSHU1kM
KmYHYBIlAujDP2xrZOpH5DauJZgsYGPg9IAzcxA21UOFtBMVSz6zLfnf4uyK+JyMMF0KmczO7kTv
hhi32oVqNlvT/Mc7tCcNG0wUbc6ZiHRkLy0nvKlvHwd3ioh+VApgCcnkQ27P2/o77wGa7Z3+c+mz
PIyV01h9avI8Li8eR5EzQB+jqlcxscAbx+M7p0ZW8f3KdVjvGN4oFjIxmUVNPTKns+mUo/yXcwqi
fv1TOGZV9KR1FPCbq4QcZIDRFeD6JRJ7w/rq5KAcIFHGDhlyWBbMOrKR9zljmTRAyPaHqjYPwsGb
MPA/J+x2FDVrpQdlmP1ztkLr8KtfLLq3cf7EjtU+eJBajYEASmia/ij6W+nITowaoOiRHquzZ3Ps
yZWQmn5t/6XDnWtuSvcoODoFLjhK2llSFqbXSIUvEXHq9MTbOYmvOxksnm50JaBe+S2+vUCXdtzl
KZqcnJPDyMm0wCZKptPWBGUne24iXWGlet/Il2oG4KMhCA7YyVYH5tGQwJpY1tIB+leS7vIBNkps
RQPETKZsGbC9ds7Z40DJ2SsMXkDgSGXh4wPh2NrWVoWHRMFWngNapiQkIADU/zezvlMKZ09yybzi
vpugI8FBNXhXK/v7eeb/5fdh0ojopiT0Okj/GP6IVmQWGqaxE0A8h8aBJmssmNpkAkzX4kO0UniV
XSdgAkJ9cW6k1dpppH+hIR+mLgLWriIhX55REyo+NcRFQh9x+JYxkSfY2jsnKyQEAZytnJPwezud
MeXiW3i6SWUKUADrVwnLnB/sQg3FeE9Kt9uPtr9ofltW7GH3omuLQFz0b0kE/cyT27Kd5KjV1klj
u5QxTeiM3pfZewBdz2gKBP++6PrKf82QLWGMAENByozS9EEk1r7Z1DUBn80/d8ZcKK+VeUgtdEK4
o0PfIyMPI2geYSDyXh+Po41TchAM75jDpUpF4/271iNs3hMHhLhR+gKGSFKA6eQLD8n/XrcWC0t5
oIpRugdBHHRsPKlB/UC0U2wfXjqQWZhVuqMKf9VKO6JzutbBWspt68ZIj5EIqZj68FrbFtENn6nQ
EgcHbGzJ+U+fVSL57EeXDjglDBuCgtcaAqa1nbYmsZDP96Lzq5fS7sCMFHS3YZ0R/WAmuEN4NwKd
7elyCrHk1QDF2ivfAXpOhpXuhEMi/kUi0/UUBGJ7vgf/N7FVp5JHVp2EyHHnCbtzu8PiFnr74XBD
/9lXKtwodvXsLQwGZH9pNZYA4DUEP02ctqFVtPMfSPH1LJM45RvwmOME/C73jdDl3Yt9pwqzdO43
IMHiwwapPJ/BXNCx/SjlqRf/GHNKJpdHh/F+2eqos/ZWUutR+fcfdIi030xoRqJeo11dOAKMUu4Q
qUaXG9hSeqx3NHxb3zLSeFpDJ94RSY+T+0X0bXQuBu1/1NLXi7OTqkMpuOy56XCFmJjpjTkhOaQN
Noefbg9OOdFuYWu9fdfMK7DarlzSvkLt2i0Fs1ydB7BqB04W7M2bRk6UX11fmu4bB3Z4IYZmnHS8
kYdymqwd2rRtN9rUiCNR7iSu3CIB/DINExQpV7CpIioJd2aA5kciK7YYJv2UlrTA3qUcWr9Segyk
SLYhx9lRNK82Rq4gNQC+0F2MX3YIRpWmMMHT0ho5Kt5723c2wsq6kUIP9fH7mDyN8W8xFlI/3J/f
rnBwszZtU3zseyFvI6S/uCy3cCVHM3vVXFvLbaRaJ/3X8P9lDYoJi4528VWKTlzBh4C0lUmdu+ls
tomZvHuHV/wqCMx9oVBT+Dy77ALFsTCqE7E+1Nkncx7Nrcs2X4SIgnMt4giZ3wEVrPR/kerk2kHC
+MjBPX3DaFHXdknRUsL5bf5owFc1FhVhQDV0gCWSpErcarz6kB6jkzoJ2UnUWLJvKc9Xzh+rQFhn
nHjojP9IZBHau+Fj5F/gRJ6neU9dvxg9T0meTn55Af78/fHEBiPJoTm7jbUK/5/4D+T91GsjeWAp
EuvFKyE7V/lT6ELEk+UB2p45f6IKbov6pAAFX0Mnf0xOg7eht4cQS/kGQK2Jy23ACPftRQ8QejYO
SELSE+p1v0Md5gC6oGoocFZ5GMswwen+d0SReVIsvBSyuH6fhPiifCmZSPIpngY726BBcGXT/1yJ
+Zm4y6jPXhSfx/ZVnO6BnL4aFYrTYNxmOF4wTufUMoHoWZuDPoINxLMgpnVBUyqBOU2jdwW/LFWP
yyDZKjFI8NQ2tTDGW84dM948M2gYEu2ZJdL0/AEUeHIF6j6mIF735Fce3wKwNzCT4feJdEAc36q1
yJ82erxC6UidgF0tWRvqDGNSzGZMPbhSFv082K9w6So7Yp1Fk8r35GEbWQqavTZ5pQNSNhim1XXR
mw7qcUEricbhd2+tL+7iZ/mpqfNpE/RI9V9mTmpKUxb84M4kMCkvQgACDYFXm97da/0bJSwtGnaJ
aXKi4kHjwSoNH7PEK1IOGMWjoGsTDyukL4IK3rYZeFVcIG8z8jh0YgkMb9fueUdflUhiPPFzJSQG
Lrp2TtyHpoJnHGCbJOdjysLalneS9n82FM4cxsdm5iQjkSrFWlle5WPpnxLlOe5VNj89twyV7gCE
4YIHveYCxhFJ1zimKq+B5QZ7+8wVvQkkbMFAXxxfoWlWtpYq0bS2hetn/2t+tuaAmHWq2/JaH/C/
Ilj5uEct2DiEugstY8mBXnCtn26gS4tf0UqW7umZrnm1yYrYIA+w75IdXLOVUWV9m5wzhDvdtdwz
OvfZSftlmEfXpEONxEPRl9dX54f9hFxpKNUUTWAwm4XIE3YznI0ww1Qxn8WlZDblPG9QwwB0qxZA
GmJ+ryuGwXli6B3pMWUX8buMINFAoi4X/diz6KuhdODdguMeMJztdfF9KWS+FqD/4ogcxXw3un6b
2FAQqJ16vKig06ucCzG8j9UyWyuMZJeV5nAaD7OWhrSg/p+ZoLaESN0xputi9rNLxsPH2llu6WxF
MbTszgi4frDqheZ/A/qWr7Fw5DJQGTZnOYlNA4UfCbQTLg4Y6/pFyXllPSO21k7bUeabvdKkdjXo
jGGwOMokSDC7rSzug4zpO7AwA2B4yijBqCaPmoYPW1Zoob50aouKjKO1fn+btzfAzPPrksOi7Cwz
kCb4V33K3G2mhIM50zRUK0xQFxQfST42ddPMhc8yOQ5sf9hg/fryfnthCBFouK+cE0muJglMqNmI
wy98858KRWvrdznQQ0NtUKMMZ22PC449JopgXeKt0W67XpZ+1Ow+dw21CaOuL8eoQN+tfc09E+80
UhYdWYIH19Ja+ft1Igd1p0qlhvM9iLUmnK00Do0x5PXW2XvmboEkeW3kOX7pbTuDX1hio0u0RVLt
UIfKBmzbMLuuBblg4lsl+KZYl+tP0WzKvpFaW/zz1Xlk1ozfWkQ0tC9DwhggZ52/rR8aAyrG391D
Ee14JSAFWbnPRRG3kq7wSqg2Wzh549yQpgFGZkPL/0uewvrjlgTMXXcpWlOnSNE5sYyGB/mq3AE7
I7d5CqYzlzL5/XE8MbE9qxMGdME53qdifT/3Ughe9HE6Hh5y+busl0vkOPXTBthvfMqLMN80fZEx
S/lSC982efh2o3P3gL7NI+0wpqosckcHqXHZ2MizZC4WIlN4vdCl0TEdeJaq+Zp+UyVi4jOIuL1J
Q1zYBYUQ37hyRN5aron0rQxqxUYKaH1TmlgmMZta5foh3M5JfQjiWQgepoTBnRsvsMJBwXhxkpJK
WPpGkkwhUsW+PlX0N4UeFnlXjG//lO8gM2dz6yXbhupl+2k53Nz645PK8990hdEa/BuIz2/rgFK9
I68R9jILNyf/+AsCxrCIUjAt79o+btg8itnQfvvMSbAKn3Za9cdWUmVmapriKvjBHSxa+9DO2Jo3
8npmk6L4D0bFahDcEg/P3AYpzhezNTX5AsveFmRVGHp/V0Zu39OA5wfdGZ70gH7aiwC4aqkG6bEc
2t8DMJRxo00KDzp6d1BEF/e6+nVoiq0CrzAQDxYAKYuoKc+F1lEcLkLrXlVHCF0NlNQU+ZHSx/l3
htJGxE64iPuQJnmiPCy93xphEEN1C/jcWp0zUsgJ5G+hTLe7zfJCFucyNXshswK8pxhNh/UQZheB
lgUCs/DyrJFIQ+lYYEnd0cV93hhWtKmPmVSiM/yY490NJmGkjUrw9OOBZiZfcXO8BdbuMSlqzWxQ
lC4TeUhP1RDqREi28tzZaVkuISGMIO3TqzctJmDea/9RHdWFbxyH4FGIwPWPDLKrVl3/OAjJMZ4k
KKQVHShm6lB1uXLrL7QejMcxjU4SbeUNwioUG/qYcv6lL9n7uzJurb9gem+SL8mzjXpaPNK290sP
HPeld6JDq1mc9V8mXhzecFX+o/jkudhTl/8Ze6jmhGU35wArTii7tSK8SjF584NbH9ruKR/hIuWP
13U25+p62t9pMjcWmqgpjBNcLT2MoUR5xt/uWUeY6Qia6G3InxeYkSsN27CyytZvUhvy+8YzzQGr
ZPdP/CxZRHXdd5ID/j9zLpyi/ctNbU3nRFdic3pYj6jUrs3U8KKOT+mB5RB3pTd8Wlbqvk9DXL2P
0H5yr0cYjB3X8oDi7EeO9T5vMRAb0KH+7uYE5E+sCL7A2AWjSroWD+D4l59uhtE7mnaQ/+H7ujKB
d4byIfSZAImX+SrjKELtSKmU/4i8cZSptm8nUSuI4/216jbzj7t85J+BM421lLMo/eMl4od6tfQd
PNvbd2oMB9iMmqRYiNw4DJOyD0lRRUpvIgK+ZAJu1+nVBi1b/im1HIEUSxVkGkM187XLwKw8VGkz
asgieaKQSXkc1pV7RrHp1IBMPpuivFDxPSgVQyL0uGCWVenDJYq1b8oNtnYnDVP464WA8FcAXqjb
SjHFWPLLKgW0s3tlMpBGL4mYxvcguyBwdxyJJBR8PC87KypcSsbs0aq7T+V23ZQ5OdqAEmFvBoxW
gWOvPV32f5Itu3EYmoCT+qVoAh2bGADymq+IxZA5PA1c7sqMZ+LpV7Y4Tj03PypHCNbXOjDnBonJ
Peh2f8v6eNIduLCQMw7gpe0DyyKQI3uKcnWSiGZURfjxDFjg/NYr93BrlT6WghAfe4qD21872WrH
IuSxn209fkP1f/M+OjRjgYmQ0zOzdRLc/PJ+e5tRx0x20r44XAjypiAKwNXumbrn4zsr+1geAVsJ
pjtk0aTt77w7LsWbPgP7idQxicaM2aNNvGWElrPoKadUoolQkcSWK5lBx2Iq3RNo7/7Tpbs+m0t/
F3Gp4J0IEGaB8yG0uMk6ASwChzI7bdsne0n1vxqEEDfwpF6RPh7eZHxWcqWXpm5rKnIxQJqU71oy
s1arvDEKkudQsVSGxrgmUG603SvVM84MMCMHIwpgKuFDdhHL1HRTGAd5Qq2KQKPTVpa72dY3zaGn
6mDbpPP9EWABwUW/OpRswquz60hGVBsdgNLcFP/0COurFz8WVgJihtrn9cq9CZdLM4esE2aOblUb
JjGIZcxKBjuHawxmP8v430wxcSH7UIQPU2uAz7kVxJNRhVENSt07RvpM5ztv2nV98a2Q5IhBzey+
ywy4VL44VeKDpcNhzV/9AYSicww4TQ2JdnLFJi5/qLxbH4fHcxaDaCgKyhlxB2baz90fj95v9Ona
Vtg+l5d7W0Q/2LuYkjBtFtyV1edKZdyCPEe/CpPghEuF5K4sBQWgEnjr8LM8uB4ZJyz+g9S+FFpa
Cvu/q5+g8kByl8MT2fd3er+POzZvLhvUbVhX+a+8hp09CDPqgUCxIg7vmh3ytQgLFuS0yDEOpUpg
iZwvhEacHNWCGet4u3GK2ZwTupziAAb8EcbvIz7sJkvFr4r3r4lboaZo+fatKmzwm20vaWx7mmMa
89RPl+cvRQ9DGkVxGIOWGDjRkFJ5RP7RbEyQ2y/QeNVr63KDaNdvNcw1Cl4tjWooUp0K3QmFR+Mb
Yq57w5sWcQ78lO0sM/8JyQykinMAw7Vf9sGRxqGF0rDF0Fte4KPcjwa0W4kCpSgcIOd6nmcORLhh
M9Oef/vleR7mUmajcGpGDRokFuNUgz6SqIJly5aB9d5u5ncfN2XVlA3T3zQwmE5VEchzhDcI44Pd
YgUJbmvWXCSV/sk+U9OvRLsc143WnFNE1Ozm3013EeJLv0SwWJxpv6NCzU6VKxffZvTskqDgZ5du
3VgKGme05A2MQ/iP8H3RqfAuaqr+bRpHkrKwZQl5Ic3kjeX9zNIA63uTZ3FrTR27SIkIsgevsu27
cJ+0mqktJuGayKutK6vgzTpMVtS3e9SgMo7AwRqH81Av/kw50NLjxlfM12GIOC8vykkofk3AvAsg
yM19Outeg69FEGHhC2Xl3v6ar0nYZNi9kRx0ge71mOU6MWl8mFvZ0VCLNNDa09jNOcaZ+TLlnkyy
o5ZrWDh1dcqdHTjuvCmwiuOgQ/sfRGLqE/VFa7h1NraH1MEZGufJ7Hl7ZhOiowRSv1rpcHY8t3j1
CGTPbsZoL3NajdG41cP4nK5s7WN63hPpNxOXZ848EjC97nO3st9iJYbynTSutewgxvT4+QBTvPgK
TYIL/U4LvnufLM9pDbopxwTatpNKvCiz1ohAvCr7sF1qaNyppNNjdEa+trqwvxmavb26dwsKiTxs
md9FzR2T47dXDONQ/BjJ4zqOIalCp071Q6wjAL5+op5UQ2hUp/OpVxo3+sS3ElT/QE5xQvY6IIf7
4aunama2yxVInVDBdwHcfUHI6tig2nYcANVwZi6LFyoylZaADSriJ0ApiaQj3Zd9RTRTCEYCUNNo
mSHFLAwIQIRIjnBzUb55dtPWtMftgFvBVHQwPso8JCAwYUZOl7hAzV0llOVX2fH6OlNDarWfxG5B
vztKVCADCPRUFGr8+q8wWn2V4qwZTW3m6njI74AMhi5dp1Fy9+WxgqOQdB3z9HHC97dMgtxXf5Ev
BR8spTJyp08V2GosKBJpcs05aOx4fzVP6Iyl5DnzrjuiFHnrj3bmtAtRC/dkEAh8UVFEeta9QNNh
pO0Iyv4iKjNgogiaiOMWq+WeM/x+WcEiDD7MJyhYZTnyoBILN6Ki4Nx/Hgg00o7Of0552hb5lm2B
YaAuWcTInXANCXeuhLnBblAsaXd1gInUyOMCIuPtG7Tktplj3lLH+rfkO/EyGY4c+z/ONrCqVKtr
M+fJ7d3vWqKMjbFCsq2vvdBUJeQHLkFXabm0EWLiO5nVbD6EYPVRYHcfwkKbCKSvd2tWvZ/SD9TX
VNH2bdnhrEX6BUEw2jdNeHcD1ZV5wcB5n3Gg/socwKBqOGgVtR/703T99d6Mut6EuxSdCOV381HA
B8ZBPJV8F0hMFZn+BBPQucIOyvEDIcF8vkx6uALCWYI8cazpfxgrs4C7l3tti4Vd39eaR7O8mXRo
EVhDzR0/c52RUqizJxHwnl64in2msn2GlQ7GAXWTP96QYZFRckRglTKLorPecpKgojJry3DAi5zF
D/J5WEAvtBcjwr5M3Jpp1u5v809nkGAXbLu5hIgca30+EBQMQZFof/HgdyEQsCklO9FMQy4RGyoy
GG7LA2LDrsEGUaqiIcVe6hU41gsA9WFKT9xHpJvOBJt2QSbEkryXm2RKIUxJncBj2fBf3RLKxNsO
vYvybe45fgdFzRzpu9KFvTsLPNbvsGSRtHWognFaZHEBjzBTcLLxL+hwauQQ4yzXnYTc7lzg1nVZ
zJSHDPSEPtI5QSP9OmYhmp9tzYkhPchelREZL2gPqnlI3iwwl7wDyNQDS7WmzOjTJ5I8idm7flsi
Bd0LGttPsoOcsP3sizqvRvsL9wopiSugyIRAdhV2rZ/NO/tJoT2YAcWigRmz/omz9mtDgKfvodpZ
nz1fBwq7n7j75fU7a89wfiJ+8zzhHNNxQwBCiPpiqqauNWsSSvVVrGTjQEn8SajjxiVcsypW+XMV
E+N8qRlvlM89W2gru45nIvIXQtj3q7dr5tHNYiZzxjM7exTB3W+wBqgUpnx4LJxLhP+Z05wBuYSr
zsm4HiIUvdRDcFii42a2mA+eCHvQpMxhfLAvArEyvBSfIpvwcgXrfxwNWGNacCdPsr0cCCjCLvb7
f3ISnNrzyGQql4Ja76zmpPkm3lphl8sf8TUfNrQXDWBHEnFKBenruZtMwZljF1IJ7earCN5pNC3T
z7wQtUfqO89j9SqSFQnT2hCIMJwRCKM+/cBrfnibuLi0uweMrdHblaShHh0OznOHJQtnet+sDLR+
/iyG21K9F6EYsILB4zuRmPg4DivQCduPxhC7WzLDeTDrOQGtuJKW9Y/daWlGwk13KTibyKrMcELi
Dd0ugjIK2Vd5anNjhABA9cRbyKwgdtNV6UMr/NSlHbv+slB669ugdfDHV8PQ8MO45yFEBYxZYv3d
er0WI3i9R6mEXPlSF0KhlvbwXh501++0lbb86MywQeu0qqanTDhXLR6ic6FG8/FRpJiF5d5HWnZz
1Nq63O7gkI4Hg0EdS73GDMIlaso5XymQSTc+BFi17pDqROl6hUGtlcPHa5UtBOQo4ZzDTJoOsyJz
azSiJBbd22og7aGgacAET82Id9tMN1nvqHgFzAOLPUECv7LrjsPuY6vlRqoWPh0/o6B8GjXR3N26
FcyP8WMrj90rZdhzAFJHFCZVc0rRF+jjGYfXQKEuGAwnJgd5iQ5cCUWL1/kptfqbKwHWvz+KrwDO
X2E1pSPIVf1zGa0oaKZM7dZq2JT42PslLMwqYN0ugU9BEEZf2bJkRbJ6Q9Wg9Z3FLuWA92/5LAip
5Vop4vstGmHgyxXgMJjScEID6CJ/f5Ia9LQY1MqXqzvcQYlOa92w6GTYGCl4R59uZa61dKdtbcy8
4bYChtl7T+OAw3F5Mwy7opn3RDoozgqMSEphwoAnD6VX3Z2hgOpU+6fj3bCznfSjg29vGJ6DZjly
0Xto0U2BU/nMs+/PJYi3gQ7pbK5ZVRekr25Rovo8vhDORm1I7/IB6G4tfCy3Nui+crj7KliNnElL
qu84kCGYy3OWFg4i2q5GDd+FN+yYY1JcquWkieh4YDIcQC2D+RTWHBIeGiaiPo+HPX8Oy4h/8/kg
zsh3tWnPaI/Ejfb8n338Q39KZDnOtFMpekz+zh7pv9wWN+XL2P7ve2zFhOrB2jBQUUo7CgnYX5/I
YJKA/ucWN7+urhCGYr60gb4llAkcPprLj0SMezFutGW67oZKi8NOYeXZXVxpWJL5GnBvENSTWJmR
S2pU7wazym+8LfGWwa4MLnzCfYwuEl+O8YF9mqc6QKvyJ2Il6f0mg6Nv2r6zQe5DXMRMmxp3w2pE
azIZc6L4gxA/UNwu++RdfbT8NUJEO18ud1nWC54D6JKdsrPLbku8dUHDOtq7HoxJGr39S/7YQPGf
I3FCGjHHhIADYchJVAdBn8IYFc0uqM77+lUQgftyecEPGYp6Gm29MJrioWdRfFnHQWLHj5xODzGq
aN4m2jOuMU6XQ1cQd39/OAhcpzImQgIlaKuuCCbzG0g+PBMRiT28P+edeHjT2pxc2BJjH15HdqbG
fLmVXGbeky/m/WI7woEe1OE/VCQ4MOQQzI3nVnMlvfjJtzNmzAsahWZj1u7QRBDdKpyPblc7njWm
eYQUa+DOWLErGx1rNJ7ux0Vr/tMwXAfC745fZ1xed8GUIQT5SXZHE0mjJKWD/YgWDorBuz9UfYVn
uL3BUN1RXfzttjdpfa6nrhMNqYQwL6kP4/srhr12frkKkK3QfDnCdJlvwze7cLRkVUr44cCoOh58
v/Bqs09QCu9PBVjb7PyHYb1ZrVTQI7CtEEdBjvSbJ2KWa4wWFkDavoTseYN+avm71Q3Lw1lKcQhW
a+q+jsI3Ije9LEMW28wRpigwCYyg/XwIQ+TCAU5jfNP2bBLY95p70sLQHrHQ+CGjcMh54mfOPaCo
ESc6IlPXmTeXdA9ys2G/ewMsSDiFRjo6sgoakLn4OZc+mFl9MAlxDGcobS6IbMjn1TJ0/+CMEFPj
v3aP6MwnP+Nw+sRgRcMU3UoemsflmfjVRT3QhAkeC77AHK7byK85OCq+y1KW8LpRgJkNtrvuRwZz
ZCco/5cWxplAavL5l78MO8YkNNpOJ6u7uYrufz2mi8NeWLfujwLhUeKJBM6WMNV0EKeS700Xpbqx
YvLkNv2UTgHNO7imYDx6A8ZiRjboU7lPsRgn9n1z0mZOfQ3mLX/m4Ci9y2KvHQbVockp0h489zaf
vKP4f41o7RA2yvoZ8ErGOdlIXVkc8f6N3Jvm7/EpTThq70sK5h/IsKbyY+GJDTEaT054oJUj+AkI
7CxyvZpUAEKn5Ez0VLOpooDt5dLeahRm4YiOTr5bRoT/Q0HAt4ACL0lQn8In6edb6j1QN1Hwa5aa
yKafqtsNOWbze8MJao+tqIK8vQ3MYnq1UdRjPA2gcLoxX3Seyj9kZZWSJzHalp/0mTqxrT78J6p4
E+ACQgNNz2geV4L1plrCZPdKLPKmmeRt6JCe0QkjA2/8rgWqR/IU5Q3qppY4btxUmFiyY2rmHynS
2M+twbXKsga8kOVWnJTFFBG06lRcGDJQxP5axk0lYc87FmrM4bqy2wNaukN6dcl+ECLbPoXsDmia
aRB9UrgIDIVjPmFWxfaGh7rcKOewU11uK7tauvbvASjdoIKER6YlsUQkyiXUL3Pzd7lyPf2LbQ2F
IOkbLNlUpkHCt4RZhQEjy8iil/9DXNMZoJ11IBsFZ9GP8OQg8YZNkzH/k0gWkVeWEM5JAQ5PJ83g
Ao/MRsELHBFNYuZ0U6uPM1UpioOIUGJOZIPwbr1cjp9icZ4mScneXpJau06fCYSliPWPldCTn3Ny
LM1YJIUF+NF84Y9gOUpmx8R/RkWHdFvCEAthKoO1VYZLI4NNBY8YGBXAm/pWAzyF8xrmVHBKdHmH
fKaWUsuckmf+uByMiiXWQTDKh11DMoGCooMZc6eGOkUHdXj66G3PBdQZ7ckQvxQ/pu4b3W3YBNDD
DqazTQu9QASKx5frZsYH0yVphbyjrUUmXbjJD4bOEhDzmUANN0/b42yBRp6946sLra0Rhsg2b7zs
WKePNCgnai0YIGJCvW9QK5rBYtPctgmgZy4CLSDWW+c3LMaPrw+GhkbvhGvDbhcVza2hkhD8HRTj
Jkv87QEBlZBRTsDNgP2ybNLte+O2YIF3bajtqf8kWGp5ipZr3Dwej2lIHctHANWo0iJqauPVmvQh
J7yWyaipPrMLMuWCriiS+l99klsPlMUyMkBFRkz1N1IGAf77EFb2bH1AkrVv+n7/csSy34q65YMM
bD03IMIrO8JU3BJ1Oz7pDuMr/FpSxWTq8xKtxBMV3YcqN9L0MO4S9RqYfJf5KnfKQuo3rTuSDMXQ
PzqRRgyWAfM381Q1o90tUaBbNkr2DT7Pp7Ppd1mvVFzUroHJMhuo9Aou2JuLRCftBxwBlqv/qytw
ayg+zTo3mF0IXZb48n1K3sKX1LhBM3+8qq86x8O8+lD6CyxeelvCGC0Ncb/3L+u22xxVs2DS43NP
I5a/ZBtErNJ260M7hPlybRfp+dCHB3E7ZWVBNkow7uNFzMXxdidsXSIyGJ7JOfRLGbnDiWYRt8u0
1L8pKoi9I4W7vis/9ZPJ98LdTR/4n1kUayHveQhJSGMZSRh55snaBgIdLjsBgjsFFSYlWG4lQX/h
EWG+JBGyRs5U3+KZMVjrkZ0NktKFKlrJjy53f2WMChSNpI6BNT7bnchAz45tdA75xHaOX5GcowY5
LyX58Dr1VwwoI0B/F/Oxjy+vfpa9K/8BCOfbYd3tSvTYGAYonqqp9mPeWlxLgoYc9WbLhx7MjzYZ
oTZl7IgOvEo1e5+G5BoklAU6tgSHFNOD+SMjMzh5WhjJfxL1kmH1j8WqPOCKLk8aL+x/TRl/TqyT
WUQ49RTa377ob5amdnRYr7L7YWojiIRS7+Y2YolIJnTe8fMPjbz+G9Bv5MCNFcNUWbT9VVteCP2R
RxrY09v5xDrw1umOaPDjeVsdxmFywK3tatDPWi8fLd8szaI28HudjpIcJe5XuzAmb2xxC/4GgShS
YAeBTJLjWnCURXxx3oXKotZgWQ1mRCMi5zsUdLGKIWkCSaWDd+DSU9VCO/PV/nZWZz8bFwLT/jpi
4VkleXn4Y9yLREVn/XxCqlntRxu0lez7greytCipYqYdJbNC9fKD48N1zv91pVbml7jSN5JS6ZhV
AwGnVi+6U44rLYB7vV1ZLlfqkBokzlN648lp5ZHhGbP8n0npE4pXu9as7c+KfhGzdFufIx27O1Wm
aiykDtDPh+tVWB0/VXK7QH0gNek5S+WwNGBdUciVvlLbwM5cpquogRJe51Y6lHf/G9K6ArKG9h1p
TWVahC+zUS7Vl1R3PBmnA+Zo5J1P02ypkifI7PuxMsLIJIUBqwet/IbDCTNpKa8Jt0zmeqhsq50J
6lThdQa7buHK5cBo9RHhbmYDCgVluutCrdhEmvybZKYnyXD2cP2S6dUwtoijReYovOursgpECB1g
bAwgNNujtzATTVFY7N1PelB3XLJJMRlWXCjsebR60M+u2Lb9b9BaHKf7UOlL4q/m+0f9wf29b/UT
LK0tZ5ZyweiK/XlNkfKqT2frpK0b5c8A7Lqc4Ryn3rvBjnXxlL/2XTf/KwxPvQ0lm9moKqgF+9BC
ng11T4G+8/L2bRoOMIe5vBKMCcqh/X7LbRq3UJgpqRB4eaTC4Udibne8/Y3pqexCX2lELppcknqA
HHVuKBS2LsQqJrbR8PSJ0+vMaE52ZQmRvXLNtNbqcoagfDwuUSMxQ4OdMKRuycUjb9scM5piM4lv
e6G2zC4uFonpy/tySRMjcnEJxVH0HN0sspcF1U1twycFSryc9I8vYLXBG/rfW6Q9Hccjy9xWq4B2
FJOd75wOElmzYz3+vPj3kxMp7pnqVDpCLWurwX6tdTvFGXRDqWmH63uHmVzFOAGXaBRsAlb/BeZ6
9PBHquuNcl+TfH72cfo0HSMpiOaZhDC6P7qSqnaiFQL4S4X6sIOSGtdJxTulnT51yk0tkJswoXii
GGaFGrfdQ84siqTkBi7oTME6EwqqpX9bmdS7/PPQMnrbx2bgxh4USrEluEksD+9yghMTM8gft55d
qaWqLQXlKFnDOgvGzRcdrwKyxnkaQhzfOJRSXDL+g+OP6+BTBwhbgv1yq7j5OdzO7hu6dNj+b8BZ
tIvZgPrjsXg51pUkk9eiLno+t48E9xa3caklEXvnN0k9D3Imah0F64YK13+VZT8fMqxYK+taXofs
Fo3I3b9kYoR+gIqS1AJ2DNzT3zACoTI9EmT/jvsOE4jL+gWIQSC44yuYwbXmSta9WC8PTruo5KuP
Rt3eIGRdUTdPpVhhu4KWMMeYbigsbk8+aDx+OAPQ2/BReUrp1d18inV4wMs5umAavcG/n3GUE0E5
xjB0+Y8CATCsRCx1AyAx4V4+jAFbezuXQ6F7rWLZPHaatz80GGO13tVkCRxzZjz49tBhbgFyMULm
fNckz67ig8PnYNoxlQYz7sVXP+dN7wFtgiksMqQaHiwEsH/5sjIX5lEbYuppqTLz7DKwy4o0bJqa
0o4PvX6gkJAgiq3EqDFUseawoOdtv2z2j1gD5ZcIqcPlXwUn8gdHqYtJ49PZBZW79dy4BG8HDrAm
ti0+Bjzkk4daEKa2Uj8YKTkiMW/HBPMDPW4zXLPeiESwQ/hdRigXboLPFnRk1n7hAcU4BmfCJf23
sPqmGC/IF1wg7s1sI04HbFMpyBD08MLYESQb8Uh0MbqXlqwjrHGKxm0W+io+DNvm9kSAs6RnfbHm
SOu0ZjVnVVLwom4TV4fkORRneYnN/H7qmQzsyt1KgFOREEF5H7iQ4+x5ihJ15S/yX/iWeSnY50Dy
kYU6BlJVBLR97w6geaCQhAGNAkfq39W0KUeqtW2+5/scED6ZvCDWOQHD2H//vp+pfzqTlRuDBhuK
zgd+GuIQhCpE6cByqY2GKr/bbo0q4XyW8cqGxfNA19BKjzdkOIHRkj6ZZONFwCuQwPQ5/VwsqkfX
OHGA7D5F/1uDLedNzt2LiqbxHfxIFyt1zSFQBctTG65SWF4qMMwCfeCJNkwUttVR/H+9yrgrj9S8
eAdGRuxvIOLcqO6YEx6PQnxvJFrySq6ztlEYS673kBJO1uBtBZaf3DeUeu9EpbH/mQEpTsLja3dO
iv/2b2l6gCdrgDKrsIwF7l7lhWPFPes0ZzhsSK852gR7gOXyRKvzg4hXq9dA6dRwtsmMH7VBp9h1
tUwQsvRpjnT/NKgjrxmt0v0vyTTZvU0dAKm9nKZmsSrcpJEkvpXHa4T5mGaxzf1HmOGRltro4bRZ
zVGvT8F3hrhJGFeL6GG7/PwnXi5FV/3CtRDpoqJx1YxaMbsWNkf9r8qSN9qiotR67h6kBbMNNvKI
R2vDWo6R9qRLXtP+3b9MKWxqK2QjD/+eqC6Y/Mb8idVJzN9yhHbJBZ1lbjTNnZJr8g9tI8+O7wRW
v2QCChlCyBMwDiKANyaFzMsnkaup0nLpdtTyr0yUaMEYfkug6G2dyBrgacMTwOgYFXpSkCiYitss
9toypUZHFk/d+kAKXuCDzI+FD5lrCY42Svdo6uGUSDZI197TjODooa4h8nlc2DObr4wBnBUcJCGm
/VVKjLU7sZUs0gdQh0VbYIzelOCPhJXXFnszTZM4joGaJTpEF1RUBSG1Sjzn2jQ3hfG85x9/NYMC
W1Qu54hSoZPPHNon7B4c2vSJKhe5vNogOGq73nATs5fg2dilwtobRYT0u03+dOhkQgMZneqdglLJ
Szd0KpTVSXt1P1IbXZ7RVPrGmVGg4AB7SlL8P/gcAqe3MgvYcONQcTjuk2WnNqOeXSnCM/3d+CLX
IQCKJN4HhLQ8Qpn2azc7sUOcobJ+Fa+rEq3WQpy5RVqvMhdvpKv2WhmsSOqGSXFMMB0hmoHYTrSk
nPz7yOICevIp4zcMK9b0jwvz0UBcVIN+4wQWudKM2USaWwtXx1jDNI3ULlpCIiVDQARpaZ+RdiXC
S8f4sUAR5VMIX//IZKwwDBJnGAoohJtFQVfN1DAKD4B5a5BXFYztI2XpwPq32CHmxJVaU/6BRTEB
eMLDnrEGzHNVrQ1hY3o+kDQDMpemoeJxPeMJeN74r7Xvl9g/irgZ55rUTcQULoiMQPiUtJ3B1Hv8
fhceeB+pIiecqIQ0tHtg7TAG9mDeLNFbcKk+KBYVQrL/ciWDk+mDykkmlMwIm+HbhNHGzflpWPUh
c+lApiSBSXXP87/kRRtntx4KoTz9il6/AKZVo4II9Jwr1C5d9hyBqy6EtWLE2m/BBScdbMD+T+I/
P8WRs/jGDRkkOJzxXdLL8o0G7oha71fwQJwuBq5olot4yFAD1M5J76KDF5kIL8LYkgHqJrVuagKl
loRPPtYJRRZzOLqupTiroJyRTAXjhPzCptLWrGGjoOmDP1PHfQSxlLlbEQTZWsCj0yi+fTdoQJ6u
IcYjCMjs0PNISv3bAD9jM/GCpuj3IoZYIVoMHkYXaS4LVYC4iGxPo2NJLbf6Uei/RgISKHoRsxuW
6aOv14BehDCH0BblEJsQ/y2FCNziUEXSYB4ycHJhQpu6S1BGLo1mlQG1PmmCwIHRcwGsJwYg2RB7
WFRU1/iirBfZ0PTIDt7yJwXd9lbhvbAy0xTAnSIOev6fMLVqYRVUPPJw3q4i/O9ZiJubHa7gzGST
ncCn+Ut7gK40flZUzALIC7wd0becKM1KZpKS+76P9jvmEDEZykjfrn52EWTqI1VUUM1OMiWrTOU/
7Ef+nL8uUIyX1ovNnbb5H/gVfTAOD9Ca41708VhL0Xq1ftGXaeZQZ1TLpJPUVtEvyAAow56wa2FX
8fwIMGNoMEfbyi1an/FGRvU1foWKqFWSqWnpdQZODR5ZQva+3zM+N79vs44j5ntutj74NTc7VT6w
M3bzH8ROyNrnWq6HHOm3tscLDuQvAOxS1Dtq+NM79a+DdeM2ezNaDTaZmGFQPeiMJ+QYKNr8v1e/
lmDGAtUOcxnJifvRqLIGNcKXTxwcsihfQjwwI2kqDhNy338xAyMtmyEtWck9ixaN1E/GtImeL4dM
f5Jak0l37g0dbXwyXyOtNBpiNId+WdpV0dfDSGJFw/fZ3WKIYzJfoNGFoYNnQE5QI85D6S4mZz1o
uwIQC5JSzcBx8Bd1mpyKfh0+vjPcLUtxw5PV0Q0uqMPQAceOgOIIJKcyFahZFaFBlM1LEWEXx5pr
1/KVi9A6oH8vRgXWRTvfd7ydr3NEXTQ0LT2J3zOb3aXfoKuh2b3kzRUDDqL/PrSOF0R0UIZRzcYj
hJrJEmGXm9Tsx0VQuDCw//JuGbldnVkJI9O+FZOS5vagmDlC0UQdNd5M11scooLgowTzDiSmXwti
b8JIgdNkG6pEswvItHOjTZWoWPfvJ+t53ZK9nL2zR0naKWRdFS/FyggVhcJ1aL8b2i5fXhTtuENu
7oclOkeBmpDLoa15BKd/i0Kd+q4L09Iu7YAzNkbaLkyg/2cej3TZYK3mn6e8XakJwjIsIJNfSJM0
LAw4ZC4e4M9fkTMNBmgepPCsR4ZLG+5heINmkhItSukeVruViV7JeaHQYq0XXGmzskQUouGp9jg4
KUF4wmTFC3dC7kr+9ezDNYUCZ3lgtgZXsDBdOUai/G4nBr6R0pmf5UB+NpVkTI2Rd1Xl52K5lAqn
IAn6Qr1lkwQhalkdtQ5f4W9f6JEDL5ph+mStVvPCzi/UxvSfJ9BzaD8ygqK/gKZ+bbhgCuM3OhG0
oy0H1gQhqJLXVhLuwHdl4H4PCJWdMS3frWmPYK2sfz30oI1zsrSF9NJih3aBGAqndc3fHWI7RNub
BaPFMMFtq34Dun3jvx35fxehh+A2ygFFw47+27OmXqxFwEJkuNXBNTFDhJslXSmXoxs5AhuMOiKg
GXXvQjrAojQYa8nVFkB/ytHcYNKmV86urPa+UDcfPoGbqsi4aTfVEgDwFlV+99uMlQVzMkbXnt2o
LXRMIc2aOxb7jqxR4Bd7Ws8lFfrADG9kjxizizwxqLb7LEFSX+RswwtbB4L9rR1PxYmna3jI6e9P
jmwx0jSjKoseLrfMMxp2w4fHJzf49WCff7ZyEaOwDykW3vCL9W4uivpBqry/MYncpr/b0vOZgEnr
4X0XXPuU7eiL9tx57ekDAzTrTpDJxvZeB0LU9NlRhN6QV20uGo7xGxr9ILZP1gd6a72cQHYp7FRc
Ol12GWFnt2sibBEwMaZPE7dhsxtEolTkSbrV/hcbQVDrtCg1I2rdOtwfiUmKhD1fa2mi5QBoav/2
Gl3IFA77XSVtENCmpsw34JLvKF6F+irtwxd59UKubhfktfc7h3ZpiXyhba5JVCdvl9NmG5UBCaLt
UKhMTNKgzpeRD1DMULLXbflvc1JAZmkMuFvaw8FjiCjHFUburfIy0K2PPqbqZI+TvpeHT6rRKuZQ
MLjKYWAZMNGQUQYeJbPH4FQCV/KW4U6o/CINskJlDYjslATiFtn/9d4zseOTCYoITHb7EfRpWgPk
+lq0pUtWmbQnXCZujYDqCoBGV7Sf7OvUzdYSXu3Dv/k3XWLYuYIpaKO1cM9jV59/kq8pr52uXjjI
ukqQWtbGcQOj2bSF3WYvybPmII1BCAv11JuEXcx2sLjdjy+G4lt9cKSNPiz/4qAzNiZMi4IeS1d4
elo/wAT78g1lE2zyBs3hpGfOjBMo48MKrLY9RRcIavfh33mZC9b2KJhKdSACkn9H8JISjgypglbi
0X4RCjL7UNk1jQXJFxkZw0FsdD4M8PfgPRoPUUiCO23gYmEzd7SXcMcakEt5dyx0QxArsbl2g23U
Hqn9rCSOZDaCFS0nVsnd4NvakclI7zdyILYUIzytrcferUrbh0f/HWXpqjSYfpbBxe7RQByAWt+Q
/6htYBm0XF4tzZFvIBQJaFK5TE4rZrW5c5Jjx2FdEEuesbVyPZp0TiWxogYeQUMhKC6wWhjjmIrz
2at/WzfO4AxLe3ZTnRNT/NcMuy5HgF/s2b8IUQaOuov1qT0tZQ0e5+ZT6GIhy4ImDA2/oEqlEvKh
MSIV9JooQNGMh7BsjlOoqqi9jC3HhCom9E4trkMbtcGNvNyoEz/UCIHpU5305sRgjQv2gWAMTek3
IwilLvtzI6NUyOpzqsjfqDYR7P6VVtZVPBzEJuNhp1kh5PyRMrJ9Qyvf8smfSeVJBilkp0qeCddo
5/UCcLzQ0LNl2Q4v791lPvP8Zo9LkBm/UaWZj94EYfls641wrQ1e/wqX5yfNSkOHvlmt/owof5/i
TKVq6AS6KSEOQLDB6dWUrZydCcjP7pG+lWg9I23HnByOL9TvuRsSx4RAT+RGPAg2lDTXcasHy7Ao
wNwwxvSGPUvcCUeOEAQIonI7UBdNNZIDViupvqeOM3dJ2rSWWbKMJ6B7eODLWpA/RfMJ4+KOIJLU
qVf7wkvDFXg2AqP1w6roebIw6PszoSsTKnTI4GPHSGSBn83gXASNtKKLJmH5/aaNgn4jKIkL4Y8a
J6EAFK/J/8UaTK2h33EgYplHoFgQ84O7f41ITxvmp3TfhnOuB8EgGIy/6pjMfeZUkh/j6fYuvCV1
AF1MyyZlfunKxwxQ5PQBO2ez1wqGewSAfjesGjEZEp1+oQyt3ufIVUfkF2rXBpRkTEhUhMBZLjbP
vWvNTnfIs7j6glZgUiet+/0oZvS0W8W2pVxrGHHipICYYE4+7q932TUiOozLkxMa9SvxPnhwryKt
F5oaSOb/GWx9uiYuFmFjX085Dkz8oYkFzFSC7yhkbmc7loS5G+/AkD1lo6Ho8JJseHzNKHfFq2X9
rrNC/5RQhoKQ8ZtPJCx/NXTlTnHw6IQLgp8XXTJSngXIgQU0HzZJNrnqJbw2aENoo8/kRsoO6mYc
EiPU+4GqBiMB0W0HdQdrzn4O715suSBMQgQxD2ksRUV6XjUuvbUL3NgZ7l31MEON+e3VuJxy5rW4
I7866qaZ/Ck6h0umItfv1OrxCpk30lCQtiAVczcO53NeHw3kyA24fhLDMSFFc76q8MhJC0taqhgX
E0NxUIb4Is7P5K6gWTUBYq1GS9LeD/TK8brJQ+BJZx7UvZb3b6v0Yw5z/jmpGvjxIaOJ8WyM/K6q
ubWkSNjEhErlNiRffUcclIBTuq7rnRinu1El1+LhVEtAnw1OG/YP7M7xu+2b2Gj+DAXqhk2ZwnIt
xz85UJN0W8zb17ZYx2xS27na8EbByEKnp39DH7n9kXkM5A75O1rHWKY9DJZW5uBLUt7EiLAz+liP
Gyfr4EITU5ggO1u0c7duhz/ipVQzClBnLn51xvdhjFnvtJA1zGwaT5xnWTUy2ic3To/WQSd35p5R
nXThQPGFr4UjyBzSz7qHEoA858eippSKCnhjwpHQ+9jYSLx2LMlKlC9vAZh3lfmGOQ/4xEIfaSBB
owks2p4mLtcspZw0UF+FmM+TMuM4nUIBB2YIoj4f1Qw2ZNB5YosSsWdq50NCp2sZqf8JxTkWai6p
yezNP3vQ3Zcbr2JKmJV9CLTNWTBpgnDVkpgH4GQc9Pvhc22PN+V2ADsmSsCxlWcUoBG1RjWXK1Ag
aCPTNmyqasvPwN4rRfVbSlebU2VMQ0Iqd2iYsiDEImFBNBHayQFsxs9vZNdGTavl6zhL9SSlI1FD
fhYp2+hAxOV416GYO9yRbxVQ2Eh1BXu/kxAkaUhlYvdEspGotN6/8CvGrwvJTcmxDA4VqBICZwv9
l8heqESCu7mlSsYLHR7XDR9brz6V9dTxMoNtxcBIyNN0iu+D+9RQ61JCECyLjHzYpenfqXJ7bnim
GkDnOWLz74/NKoUONkdyZWrDKMBpU1+nEJaQkdnjTEPbrSqN42av/vKJGoOrWdO4+a+Ee2LTkLeT
Y/l+eOG5ChnooBGsuKeF1WohGuQ4HDMQRF+95lTrgiXEaTaw/6YdYA/+QsSSIdNDHCfzmMtn3S5k
5AeFBdbya2JlFK6WvwRaG/tLxecbQfcB3/7wOs9j7Qy6Yq1QmTROggRxVr8lu4AGQh4gdx/acQ5d
IJk8eIjV8AJTn/yIqnrXdkC/SMaSU4tEIAqGk7nUp/ACVhnh6KtmvAdyqEVSMfCo9PxHRHn3ForG
wMKNe3BXo4oOPr4pjlRg/rgKUJwdNrW+ogsE8YNWBwc62ucYjDxX4dkXakach6LSifMxWaGIxuEA
xjMTooVWNY0i5D3yJMFgM/1SLdxJruSxMJCWLVAIH5S8JvRyxTUtS1F3qWH7iXHY6voaztoa2Rvt
uQ1eV5z3Yat+xtXMbGqDx5pY1hopwEfvBOVS7MB7lxKhC7QF+IXX2EtKDEDgls99vqURxUPds99H
rqW2gOKfV4cdYYdbP4iaYp09bBgbAfeFTsEidCe9WAwxJWA+RobuRyg8JULu83P9pePKutEtsEt4
6DsANxSwL4OaV70RGJGbH3k/3nzaUCxY/kJfC8+jSo88JRoimcqB5698g+MH5A//mYAEOCBOCqlh
StF5w2g2ytott3yuFe1L7a7SgGPF66nrPY5LBKHAZerQAK0oB+dW+/5lBfxapRv696R6jPHAQ5Vn
mN+v72mKgxRCp/6rFgH9sw7lzzl8bdsMWvOwCX+zHWjtRQgAGM54jx9w7SfQriUiuHUWWppQBPML
IZUVFhcncIRRUtCbVZsckaMPoPEZeGnQYyz945NdfLAYQY2719nVqX+z0Mv3lZ37frDw0BxSr4ck
FM6mqpRRaSMFOZyhEEFl3KE2ZC3Ld4SDL/cITS05MPaE+y2DQLSnu6CtLF0rwVLvpxfyUDvQ8uaB
y7r6nGwxEYR5Fk9B3t/snKwClckx09IKylDmbS+5Cm50ZKcunZAO/l+92jGsPPuRGZI07edYjn1J
aq8qZo38OwIX2X3SVS3wQ3WW/5irIkGqXth8cn35GiUMlQXFCBvsl/Ti3EBhyVBZJrbgP56RR6BF
DV0Um4iLlG7G96dVOy/nlym7aOcgyYMq2zW0ttowrddRx2q9Bj3fpMNw1KVKzrgcyduFcIqVBHEX
bSN7QLOoaoW2PvNyMTD+bIlPLZiQtRd5t7oqmXWf3wUWLUaHaZvu9mfC1bB4TH8C26XurNJ17Ide
4HmRaAMLExTLUpGAz5KyH5JG4eTlPwngtGdb1y8dqo9C4pBiQAKERt9EDbg3ctDlwISMrQg4idn9
7zEJ73dGX70B0N8kLab7Uy+tXSClynz4/7yeXt0QMi2OlSOIK1s88B2U8jl5IITG1ONd4y40RyRQ
dYzsOiT8MR5L7e+DHU1PfTZtoFqg5C6uAAYOV2PvlZ2PlkNmWXeux3jiRH8ORfAtuH16QGmFYrJU
7yR3MxHU+a7AFlXlgfTbDtaIJ2Rgq21FH+12xIYTylIxnUDfMqcQXzPDM5hD5s4S3KLLB3ey/8B2
yaQljzJz7kekgcXOV/dNiM0eK1+Xjl9+JYcS97zmvF2VV3jRHCpIb1AAEd17JI4Ddre3C2lsXYst
nJKVlzR6lY9sRol8v/s7DiJhuw6LzfRCZFR8+XDKpte++J0XntxSa0ydWkqu6rupXJhfMYIDNGc/
IEkztby7ohtqN48g25OxX2z+HKMtfeoE77bmlJTP6WdkuCIII2sTaE0fx1exeY8cicNBKaTpfa/t
p7bXt0JIAXCBD2P/PObD63TaYNnT9NH0l4X+KzOsUo+BzQ3OY/NCWiA/xDHe7dFZceQ2wFJ47y+4
Vn4w5o8Bd1KWeUFSyYM3te4p2Bsnhn3rtsrr7prpHMqvJK9WEGbY4A6hBlHpDcY8/OpevP1Pus7E
pshJdRr3h/KZQSD2i0K4uBCvX3ynTYxQ7P92RYmPwh4eFOkTG7TPlbi33FCbuYRTnMrCdjgianPF
ul3BrA1fk+R9wLBWxsJzfYj+j9YL0avsRL3uckMlMr5Vsl5cCqYrtfNQr8Ruo4G2ejNGFjgkQOhO
6WpupddxKQIOTvq8nD0SqfgP9xnB3pe7Li6HBwPf4lldm+dk++HTjDihQbMk4iiXBH8utkupli6v
lf9tZOKb4esxmfQI8Ato1j0uwCpUUiZaP+20bq70zBDVPOOtwHiERdVAF3dLJ4Y3Fitbe0Wv2iMc
P1dmKmZakAtmQWmvK9A8o+64wwVOBorV9rGnoC8Shejtezxg3ptW5e0HWFEON48glYi8kcRUQD7I
Ghrw8dfZ5DAJaMKqkqNeHUszTYZ8MsXXXnDEXj3DXj2xTUiv7DzW5pm3D25RaI4PaIOBzYi5cfP6
G7PR4U88crT4XWbOQWkUsVZ49vOSQhCg/tpubYFTo8XKkP3Ia1oZuclC+L1985Vlz0JgferutxqB
5mbDTwjWd+gLP+ciIx65M1A74RMaJJA5zzM5ciiY9r0ToFIEPiH0C+CeBiB7BVSjTJC0+a6qAwLS
51aqeOcCeixjkxYKQ1TPS/4zCtcty58EQw0Ax7noWdEwNLKxVKNuIZmLWrvgrgGCVQstlbhX9wX1
kJVa6c5StnNn6ACJIAfmmFo7GRSNDBQGfL9QRmJGGXWQV0h2nlwQXaXy/9At5V/GP0qU0iZhCQM/
6NrSMstUcHgkVyCgaKe2y0Nr8rn8LcK7MIiPMWU9MvOdS9yluKWmrFkNyN3CddM9lV5bUItIyTgA
CwfiuvnMM138vjY/DlgQlhlxpovMkZR1ZRgifcSa41ebvJu/sV/XXzfby+LSyzoF5CQM5CTRjQxn
TSDekjSnxzs30FgAvPsfc38mTqea1mc2OhgdrXPEbroa/6XD21YkPXXjXZEzgy+KAHtlojY2qbeP
0n7KXTrrUnmN03UPP7rNUl/J/7b3n83uO/zFooGPj8rV+o+sp840bPFXAuvNw/c+gB8pdk9AOEMA
Y1V7pbIT8iaPeEpQMLuP6H1zI62UGt0fBO5tZw1l5saTVQJ7axk0Zk4aYpre1ayFvwaroNkfoK8i
nTVSF7pHdcIZZSQxSwsL6cy8ICSajOI2hMe3hV4I+xKo4b6eayV0FU2Es5zyNNje7TcXSnx47ju2
WvY/BVmAx7cfYLme8Zu3JBimYm+eqbWXpxA2FCD29RSeQQSk/oPVuxguTng6XLCzN540mjRrfZhM
4vzmsQ/i9pwKKPIIOk1pB6N2XMPlZ/LganWvSD1bh5LZ9DAnBLnemTqQsBxyplVN7PLXoXv8Oph7
VeoFqzhAI09wuCKEl1fs04fIU5NOpO3Ddf8WzwW4ju4euOR1lGaY6hfVXByqudNoMVIGywZUoT5L
8p6oJsbgqo6A8QYEByGtT48i5zgN7RxZ2Npe63yMLwZyE9yZoRXyq1pKXsL+XousqtFy3xpM6vi1
Cr3Jrty+dW88OVcNzkD2CO1/5cb8raXGIY65kLUTe/6IjTuTZLJ9MCaSHirwEkD1UZfUaD/5NzQW
Jom91GXnBUxiWQyvMqX7Ado6OX9pq6NA+zvOgbTxOM6hVfluqnmFt82sEvJHTMzP9HPz9L8rhwD6
m4FxHWJ6VeDjKEu8Wk5zpbEYXO9/A8HruQ2L+xBN95TWB/xyl74vNZDx9NPUPoJeN+iVV6MAPFZy
8rTgBFuHBTpw+G69uy7YG9zOqk1HILwRjJDvKBLkZqcHfLTXGljUYpjg7WBSNxTICAGduFsbuaiK
tT/YLPzAdBdVuON2xsqzT3mA+K3+kJ13pY6jIyUIxtumYfBRjKxURgw7wVjCA7pYd7fLLvXuL7CN
9owaELKPSegeygnP0p8+2a7Y4JyULxd6439pDDpRaAnO5j9Sty1ITezvJGrTrmhRZ7Whw6B+PXqu
AQvJfWsPako/WZ6ojRMKA9Y/HgcH8bnmh0Mi8gp2zqomise+Rr0UtrNaKWVptwRJYLdk1kF91f6i
N7ySPrc4BSqDfTF0hHPxe05MoRqNHaIs7a+/tEotkhrmWeptdtF2jYiKwyb+uJW8OGnx+BIdU4K/
ouvGA5Q7PO0CSj39Z4B9iASi6OPUY5Uacw22k0yVMv+g9MqK1ApMkgjXLG8/iTuHXz7ns46AqB03
hop15gbuj0qJvVTAXSY67kwTyBY4jgxjeDoT/Wz4WKfyeCzoBjWZYpm3lrqW+5iMJqA7siPwRebE
KYEjsQHWb3/O9LrFyE1/V1VXuNYoElOQZjF/szOl+vLf0LGIKuO0Ul918wmFsqdDDw6F0q/YG1ea
dYvpVSLP/s8mWNNcY8PIv4yeArT0cjGIgKZ0n5NhTMliYa5OVQpRpBMhKZs2sdFz1MIJe3II+zlA
tzfcslEc95kO2ezNSTjpriEIgDW7NVJUJeZVvwQCECb6bfVCztaeZBJbSbakAeNPMKa3tE5Ex6S6
Nw/gkLtUvR26djACPB+9VUzB+SpqnCMWD14sflw0r8qspe92W6mxFvVqx/ysrWzk6+S2Tpahx7h/
vHkLkPB7rYcJBJLejoqyeItOAjmWlvBoV7ozw6kDLE7ugDJoYZnSJW+n9xLxP5PK0egg4XEC7a9P
elMg395NqAN0vMZS06hbBTmOU86Yz4d0IeYYgBTPCJeEM0988dJ/YQeKS3WXnxNd45wufpk7l6QA
m3voOrWBkjXwFA/cmaNeaYxpZnn0Vee1c4IxSWh7odvbog6MvC3IvbBiNLkShr4J94sw9oOFXnod
DO4Nc3tne3qSQZeDWubpToY//aePEw8VJw947ewARhLqQmcP8+nwV+W3Bgoti23EmSuyxe4QCZO+
tMlP7FpupibeuiBeKp6xiUw45tFRnUHr8jyhEFa2TwHjd7esRNVTYEYaxxCmdyuIgO6we2G3RDU3
PaSyvyt0NybWZFTqiK4Ye6XXELP1mcEPAwV+u4ArBQ5bZttqUOuENwGaWPcHArS6IxNB6Gi0aOEL
NO/a67weu3ySfQ17HkdtEs2/xLZUs+mtc7xV6uxER+sXRHXwwIVVzintBNMoK6YKxEf95oWKN/5P
1q/Sa0ehQJJDKK51NBkZFZuZMtlBIw72WsIi7wmoZA0tSRg8IOiFCDniqoMfgFLN8IONyopL04yR
9YNQKNyOuuFuR5shhDgkrRBIK/LwKsAgzLucCWKRjbhUckozl2B13RpohXo4ZPObepk61QhvDGya
U9v+mnyJz5rO94XFPjsepcNYxo4IlkjPQQQrGG2mzjPmczEvye3hTztdiVxs5b6OCeoAWkjLUjzm
Xo+0/YgJTwqxddnNokgm8x5S2adKMEyYVLXL7LA0+FSIK+aig/ERhDNx8qAauznVTDSRC8UEclUG
8XmxwfdApGzX2kvLdJDDPNOvl+Sebj4jsrzelweipLodp9GNwdNqZjVCW7eVTkTDnFF59sWqyH8C
7V+JxuJIhEShCL5Ds5Wg9Tbr2X8PPovXTb9wTytLBmowPKy5/U/h6WP63dCnaPxwITV3xVT2f0QD
7kFbz8EXTOOwzmxUQFkS6dI/YwmnL8e3p4dka34VGdm939qJDISOmhk3SlOEZXi8Ydi/sRBvJ2sv
ThR8gQSx+kDlel9CSx5xS12GFBrnm2vTSfnOK12boMZxaVSRmUf+zgytgkFGM8Ni1ptgcPziD+H7
3rhW6jeZkQa7HyC9yXbZjONCB8NG2CJGfvuiXxoASHqswDMOV8a0Gql5AVxXnumW5YgiTXDKymdz
T/a95gLlgOG4BKkkLSg95161Jfmjgd/7N6UBbnZBHu8+sI7XhTV+2MvMuSqm9CkhJLmqzjo7r5iS
Uh4ZeOxiKifnpdrxtTlAjsVeOu2A3p5QgVO/+XuShsV9AMAqG03AjQPbr8Szc2snmTfrh0SBt/bk
FnXXY95cjehGSX16nL/ZvZTUe5+hQffa3jzzVPpALoqem84qG8P9Ka/K5b5ghOIV47/NWapX23hr
GsTwe2C9P+uvV6TkKqmgvUrmrmTKRUzxIs3FEi4SnRsmc3jW7xvYcLOjRO6CwYNfUuAARCOUQH06
sHXedZVA2u6AXm5FGdZn3fVeNTRmQJ4i/fgBAiHh6Qb0Y/fzez+4v2DcqFwqvh13jJBDxF+A2HnN
cxYay/DQbpr+rL7D9TG8+7eT8z2cuqFD6VEakRROp0i/7qiuQxByGlSzNBS6GJvX7LIxGHyWtoZp
od3MNCM1ziPFj+GCKkQB/77bkhzi0igq8QgWpuP0DdrQo2tiVUp+bzaaDLt2WOzFutjvJ0Bxz0cQ
hqDyAmHlL/zGEFws6k0tJiSNtCHu1Gyw5eijklDlb9Icj7SETXrZEpt/SbPQGOy9uRxw+m2UCQKa
eKa3n3TCEStVikE730Vm/v791HA6pJt2YfZa5tlPgqwe2J6r2SNX7Zmz3xrnOoZdWeaED3jZXgIj
Kpy6fVIEN5zCiG8PYoEfslR4YeQ+E2SAUrIXcHQTYHxhu7oWyVXydXO87hz4v3RCPbfJ7fbLeDGL
QeMiO96IPbf586KWHV82VaJp0XvG6wPylqt5Ib3V5iMgXLSad/YLfBvg6371mQypkvaKBL+aUMJ4
zsCeYNgJWX1UWqMFnQ/2eDOf2wmzblz79E/vNdGQZR6FdTwnYF5LpGANXVcFF1M4VwiDRLQ1U12b
53pQYF6kqAmzmuxbhml7DJ7Uzygnu+RnDgsSCOsvGrkiUK6XSlsktsginasYVHRGqz84e1/16dmF
D++5fDiQiAZvizCkBb9j6zZ8T6oIN3QCjQVlXt6lNkWJ7RQBi9/cMJ54pNs+zZ1DL3jxwuYXurO0
qvX3i2Zl/YR3sJHcXDr4LWxJIahnVcnObuWd0I7W3lZ+LtM5l4NR3FeYcBtDS2swXS5enxm9gHl5
tKTps5tjWI3i2i7hKoPhBBOUsb5tOeSumHBKwYVpe9CtpxgX2FO8DRelbZZAm6m5vUgjQc3vAyv1
btvHWi0erxTY01OYQQW4JkJ6k2C4TkhKOZnWDtiwGoCgcgXBw9e15RXE8neZJl9BQQzo0zHU+G0x
r6gOeFbY0AVNL2h5vO5bIk2b6GrauNho72UZbj3YbMk8sABHrBiuDIxGcDeGsQ/uG3KSjugR+wm4
ceSMGyCeHKncn11CTRb4gMZKEmRFFpt+ZGj2h3red6iS1Ob4bJ8PaQSLQ6/3YoOLzvOyDHWMrpGF
6hkzZBsgceRGyaUJrOfGRRAQcPnHa4a7Lx86v7J/lSX++iDosd08//eoaA9soxKaFNcIwPcF68nB
fvSuPsNAi+kcV+qLhdZQn6pMW/SnsusMTi6mq+1HS9AhCw0et3oDw2+4jhpFglRSNEIoiUn4HsWl
K4Bl90p8hgSbPw+QpumPzdj7/TKtyRsK7qTbx2k2xGV+2xbkcNPN4oQigeN6TykKQt8qPjbdeHG5
E1V6pJ5V++48Sy0Zk+wcIeTT/s1v81Jx9LL3L+zxDiJBvYmF9NA4ZdGlWcwg2lrImub8qqxlEFBT
BSfGfkzIycFCjvPcPTfjxqjH2CLW2LFE9dsKpSGO7XLVJDfnz0ubprZbQCaR2ZpSJEG5cWTTxzLZ
vcGULDiqh8931bUSwXwMwmAm9/WtQBAoAkzbrJ4xEC7wk1fIHmNETN6eb4cokkamfUfTV3xBkFsH
6HVa9F4JrJbTcVGQIOsWM9OKe5BvnpoCdR28/HRNWp2Foyw244wNItIt3mkd/ovafO2kUhds9ErY
5OTFXXC4DCfaJ8TXFBWm4pDF6e+1BDXXb7p3/gGh3rcGQkS/TPwN6mSNGZzO7fQL2Ib+K0PpG4IP
HMtXC5weADXvxNf3UAdCmtmciov4XgpVaKX78Vm5vevhIO2cUXMOCCViN1DijNukZ4md56QUjNp1
YtBObN4zJQGzu6LoUJ7Og+RW1ElVc91K15gfcbwSQ0VuzuZ3fttkV1py6Cd7915bR1IRf7ATdOn8
D19zDo9Wc2O2XV6DWQPnelq6D550V45jsqIJuTgyzQYgobbJiZ/ujMTtGL4k69BCzgZh2IDtbGWZ
zSFI1kZ6QAcWCM/Oaw/A/KwqsWZQG69yd+4wOwmxEavCincVWkZENhtRM0gVnz9k78/S8AvWZHBw
zQZthwD8YTN+XBh4HkgW96DuCjYsB++YSHdakqbxX6Mb/vRpEPsU33T3tQuozhklfitFhIsAa7jj
Dro2xRdZC8pkypse2qODjfjbSO12g8ALxXox/eE9OqeNP9jOGv0fLW8JZFW1wMf+V8F+5RTUhPeo
KZ/lONJEo6MzJdloDpTN9dtXSvIwCjbxQODHopAOPQqjPBSFNuuQkVyrV1LDr+MQgOvvutBpTjpE
coOMQDw50J82axYgvPVRB35jDZaVlwbfSroqxe/eqx3n8ohZ/TFdj7rzhtOb4IJ5IFHQZGtNN3Qm
dk3VAwbwhiKghHrCUroUdx2gEujFXah/8ekZfFaDdDHLkMVP5Z/hZ5uMavegVTty5czcWrX3IjHF
QGMZHIctMEvKMd5jsh2M/uO8D1QevHZbJxP/9T9nPEbQvVz882cyFBPncf0BMtLHUa5V+2w6guws
lZygIf3qCxLiQ2VWvBouF+3m92l7BwC5HY+TzADD5cMpbxS421byMKSsFUacct9KYJfzH5okV10e
EmfdbE5+h0+HWGfLt6FLjSu/mCZkjXtgB3I8ki083jRlmcvdyosGVT3RuExN/A/jj7xlSvFnWp93
l0zTtIPk0aEHNvMZOsocbWyfBM5CZhsgQX5UFkddeIj6C/vHbKPoUrNhXDtH42MhyDjXcSr0PhjF
IHcd7goSCKsv9Fkhr0vMnG8b4BH9YJohC1kCyfm1JElwuW44z9Me5VfJBINfdEk+adRP3V+HCXYh
jWwdynbyMZ/BtzvW/EYuMfbO5ZYDO+0JaGHskbR1whX9e4T1j48n9wumX/uIUxdDrT/iHTpcU4eW
pMhk1KKgx/OUB/zQeIKDP7v6hWU28XRQLV7gLq/FdjsPxH2JGIVbs6OY6a6dHDFOl4IijTTWfitB
2zoj3WVCabTm65RNe0oWQD0EMZ7lEVPevWOy3H6qzUYC200mMf+MgcgMM/qEe9uRA5n+WRTiaYY5
5XpXiuo10mZKUazgscc9mUzEEn4VsdlYWob5FWHjrEeAgucs2uRsKev42ErXqmCAJ3grhXb65zhL
6A4mEKVs5qt1whOk9uWqp5N+4lhg9z1QcXyp/AeXw9yLjl43XATvTh7STW74Zeqp/cStaMtWw7cq
0hBnN6KUDp+L4hZWoRQBLKOnxtgan9IVtKdqdiUQ33kRo3RMiXBBxYXIk6DCOcDWu2Xa6oOE/nWV
aDF8wVEzKdr8v4j85HyNHOz6nJmZ52Fkaj07yotHPgtyrXQzIuxW/zSDwcmjBgxs6ejBHCH6ClSq
zVPPO5LS1EH5vaNHdZsaG9UGU2fHW5xlyd6G9EgtOS7zOLJraly3NU9/y2xjZFBPKRkbwlNSUDWW
uDOaq3tf1imdGLFPz4t34IDv1Z6ri6U7RbfhaXXK8UUR+UZxZbnVx+PPDcQk6BMa/ZTMQLBsIYTn
TpI4TeddULhDSNWjtzkMvl0NMeaQ6M7ZcyONp0dQX8Utq9lmnO7yhBsYMNHffXe1UGbg015anWC5
00kMAxd90hHW4IDvZfRPS7v/OwXRqEdedD8ZNu6TuaHz/cuDnhyPjmgFagh1E5SfY3aMi/o+iLVx
lKBjgOVLj1W2gW/Gf0r66axukDxMwESyoBaZpViRxx/EAbaC6+/bV2ExtTlOMBL2srHeuXTGxIcM
XzrMtqT+N3dZYdXXrQhaNSg7niKCY4EweJEBok/AxRnnUfs4gxJ15aQqoFaAOnH++WZoRg+Ndv9n
t6mt8u6iVWj/hFIHiGu4N4xQ/7lOWMjq6ftI4GYU2Q8Hweqr4z/grqCCvWK4f3GHvP9w8s0TO3fv
2teeDHDfxvAhQZVSvyjsKBMHZeDCnwvJKZy8DbGhYtrWH3C3aRVgAFLvQxl9W7eaFshFgjH16hD8
FQZtXx99H3BA4O0lLxuBgembjzIqKYq2lyfS5nbU6CgclfNiSX8BvkPpIWQixi2EUAPMk/5v78MS
kJgBE788QfAF6JDFj9tokeh0yTB0r84LmAiopI6IuqNEdbPaB0jd5y1ReVQXPFKkBzP2y8FDr+ny
2ZQ+bX8dxruUZyC8kESklZQEGWMPKSxU8oUzZUushgdMFDpp2nNlFOE4q3yY3Qfp8asO+JVOwwcx
85XDLfzmcQOX1ygyJ5m4E14RgKNjDdkdFwkg8gxzQmARop6Fdl1FoiZ95oAgLk1OZCgrcEv8GlOA
YEY7j/DPQLzAxiecXdMQ8cFyVyd6m3QeUV6Xw8tSAPjUBdQQYDPvYGHX45KClolMsUyvUmN2pEsu
m0c1d3VmTmDYgGZnAVbWA6J4cO+mRniehDXT4aHLs3r9lu9niIgzuF0DfgpWqTBc28f04cVvu1H6
zqLmtDsS98JwZeAPWyN7G7d8ika6RAVBGdJS25RnllZdN28kpVoKY9KS5LtDweDVvB7Z9TEIcG6P
/lYw/WP1Pm/UHbOj1yzNRG28iTPNJXYmUEeIakVvcq+FxXvlTj1ojIndoxkTI/BY6ubQMBzcetGl
Tyvd5eSo/qG5be/B7YHWlL3iyxmIR/sWVfiz7cfzqSkdHWAtOFSjpro0QZ9Gf7Z4bb8fOPTI3wPf
ZBwzVvXHiPoosRR2G8o9Wv3YE3k/FXd64uAraSJ4MhlGPlAtZ4/bPmrbZxQ94LODVDs069II4IDf
JRVss0OK0gM4HCBeFpa6i4ewOvjXM37W0wQRhPerevC6vtxZXxPcbZbfINpa2U5dfLN3jx4j8L/M
F69dki7IptlvL2SnboQvWM6y4PnBhuwrjs4xOPXfPhaqOEDpjIRInx5wCvrTkmGwfWrDfj9mXp6i
PF3bu18zUI4TERXD9bHLVJ8/XxT0VB6jlEH7TRNg6o8BdgV9DS0uJK634mkASkY1BGuU15Hji1RG
qE5R6OcdUmbfKVj+OrZXPv9bWrRcl5A3v4SFxOibBazvAB1GDSD2KAsx7eyVS4hgLeAixQ/ALly5
SK+hxMjTV5MzTHmPwoZp0EeVRriuQvPs2YR4QZnGRT+EbzP4LvlrDxLOe6j/+A9u1nkRXf4TTew0
z/BYVZqPJ6/+wuwhbgJtB+eXpavGOWUGXYXCXvBlmFaG6AEahWrnpS+u5VPacJNGgZonhjS6I6Yk
Nwcv/TG2+XSmzH/9B5xVLXwTJ/PpG9g51k2gzvQnzxcizXTApE0QSrJtuILL5W5eJ1vJBC+Xuo5V
JdFys0BRLofEpYdF/DsGGMsHpwUSCjGyJj6/xTcQqDdz+VzlvQtDXWFIXtjZRYZKLn5+jOwim6EP
XgKq4J+6Nx4RtG2PagOooJYXzY/QMsQYEi/1RUcpsd0PgUZxJwK3rsMuupOZUvK+wpbkn/tMeOl0
xHAyqCLf8reVBdrnZ16zIWJYMGhq2mi4c/bg597yK7Vu5iuLte+fRRh68gY10VUPAUITxjdGKFif
3YP1FnSiBY9mkyrvgOJhWkDyGGOk6dChGyHZ5lSxabjojqKpXDLJNF8rV/9XgWohAaod1uqDm+XX
W2HCV5Q66vacIZjPznNRxedk7ygoCifkRfS0GW9uX/hgRlW2gvXnUTRutejG/aJK8LT0/UDCy07k
nIWdjOeYeV1epvSaKKmunpo2J7FmFcRPw1Viea7rzQ6apz11RF281KgbdzlkMbu0Rp+2Fl2JBN1D
shYU1YLBefYMVopIAjn/zzpNYWvTFECzuowC9MO9ZmlZIActmsSd5Fu62BsP6YUUFM7Td7EYgtft
8iLX5s4U2ddODx+PCD5SMsIeMoBbywAZDWzc/7Ej4DxTw9yBZ5Su1j+0+fVJ+AZvsF9AVHPczTEh
aEXQLg2Y8jVVMCzPAEaY8amIyur0jigL61oqGI2GYLdxetJNPCUJGpY4QoT1v8AIDkr1ZjsGl+VP
Jv+deFtB1eTAba4Wj5rJ4xohN0PtySO1WvCb9lb61FEXC3bYZ2Rg1XUCEX00Rh5/O6uhYz7C08Fg
7al7lrFsMesSH1Lm+4U+XQAKjQhxyPgYQdYtauWmzS5sF+RzcjMq6Zqb30n4gnInHv/sYAh5S95e
2WQyNlgcbNW8A7oOHmx0xo13t1gqL1WRjswvDVsrKcE1CKFjssk6uEn4LrSCRBqlgFSiiJW8idV9
0KeO/YJXqnXTPYWiyXYeDSsRx7h49kmfuko45YmBa7CPXKzerSp4Tnq8yvCaJr0rdGqTtyYJFVBj
bqqN4XwKDluF2MUy8xNwRR0xuc3mMgksZofcDJR8MQrVXLOxGiXIsSRckPmsjeq5i+fcpYy7g4DW
Jo67cm8RVQjcIWpO61JcAd7fxlwa8082eWtwH30C3SFRU3aad3woi703Q9Am0bbzRjzog3FrSLOO
m5GTGPteH3ntqqAyhv8+t6BAC3qUd9lvY3oyOzxhAtsMmetq2Kirnc4tn1xtTHAn/Wx0PaTISlZn
CB8DfksT956rbzTjrt5uGf2OO2vxMSATfEf0aOSH7ySDWDfq9dRxbKxIYKR1jALjcWW/voK3EyRi
tRb2i3bMi2wNKyUD7BUO0WOXjtHPbY5vnj4OkcZV0COENEpJd2By1SkQeZ+80F/MLp+nzLgypL/7
0JoAwb+53NB7KqpEG0kN1prDdEqaFbjHhCDWXXROtHeI3rBnaCm/2ZoqHgKZYU7Yge9TvVIuQu7+
pn7KWuSwVP082bXTruVw6FilTAhee5ONwM0xoFgR/ggZC24NAW1tzVMJ/sWd5wOTRPu738X9RXyM
O7ZQqW/UhwnxdOH0A4jVeQevEZw5Nq+WlGljA+nQaFvA5bJwmIn1t/qzRFoDnnLZPbo7RBj/BVan
R2b4L+bkrZCpTWSTvPNXSDHvEASyt9P/hr4ChWrDY/sGTmRaOt6l7swGDPNa/8iqdJdbIIu6Ms5J
ihEteP8kwKsUphVsKxIqYIg0+87Hmzt46soYcDSFzUlmYiQDz+tt5E1Zwh9dcjYCZjVQIGJGUdBe
xus06QsfRu1yTFDGqj+9uy87+bOAIG59E9DX3Wy536Uoa3wwpY/Xv1+SYDS9ljUCfukvDcgwWmnU
0lkHb1v+CqlGOfIQFIs6xW3V/1VmH571PMvd93GMoa8YvM/2WUfVV12Nq/mYC3/OAqc75zC4wYkC
grDYwrf0YUMcL6F20W5uhcAZ/8fV/l1Oz6NeEuAHiedUzrmyF9JPCkE51/gTOTsUsVcqQgOkweIi
Xp0cVvxd/yd3MKRqAIwHWJW6SsHKqM++/OSnigLONKARz0l+1L7a53/bUhlnnrs2x7WkdUdmc/HN
MD5JjBIXnARiPnZ5ebBuJoi7u+eyikeobjm7MBl9D/D3oLBxYuL+ArxiVUTnFqP5j3EJvA7quzcG
gtdNAUoeCs5WTsF9ish6A3xgI2ljx58f078pdCLKT7TOfEh/bzAug9Y0T3/YVtaNsjHGzB+5PhYY
6yfOLclBfRrGKq3XGolURYRSmxcYjbj5RZKCRZfXwibcAa4E798tTdYNKAtHtRM+XQRu4mYcQeal
BSfq2dnfTxnBZb4Gs5GeSAq503G/9TzpRTe/InAMrz1/Zruv7dCX/bQFGNw18fhbpaulg4BeuDVL
lN2qc/fKAc6pIsX6Di8gHkHXcxoFz0m++RgrzQkMdzDPVR8n51/4qhJZ8QJe8gNm50T2v/OqndyP
cf+1Tl9vRtF7zMaHiTAoIIB4thcxZY6NAj1rUzBazW/0ghkN4ZR+o41mrjLC4WjKcL+t3ZodDAoX
yPGECtwtTUl47tKqpyHiMWOBdS+apKxbNiZwI2wSR7C+5aZosbip/7ln3XEkZ6/hzVfzkGIpT6CB
mRaBwoePr5Q3oztKNYv/rkwpa0aluyH0WZ8ZGxgi1PkRm/QuGXc08Moq0MWZM6lNvMTI7yvMA15w
qmSjt9gyuwy3kmaAI0bj2HIPrCnOJJjmYCzIIi/HsNqTYPSz8QtMbv22KF6AcVV5ALafTyRaxiEn
+qYQXT58Xf4PLkkGltKt1zd7bvrQas3grk0hgmVuJgtQBkbZK5ivRQpwRSdoUfnTLWYKwDkRIZ1c
CHSlQhv5DDgXP4Zx8/W3qM04UFqWi2onl3OP//FuMbW/1eQayYz0TvxtKNsGqyPFOWGbI4mpOUg7
Agrl+bVvSOEENsWRMMh675KrPxyi7aE4Id0OBegcdeO9PiJlElZcAyF2rky06T2WsGhMSqO6uPQa
khYmycP5nmxg3jRro4u9DUfgl6wO7SV15LO2uDuYG5CIgmgrshaBsB047/dsIoBDbWbT/68MUZ6T
izRBCcdghWRv1NgFA2Y0/cqopGd7uz3ap7FinWWwQNrNbQxL0l/a3Rd68v+YxZi4KmIY4VePkokb
wLlgOoQ6ri4PMpd68sQ/ibwmuem6hXTCJGWrGHGQSVueB/fLwsQ2UZ5Sb1bjrsGLwj+PyzsB+wiH
BmtQOpxMvFSfa1geB1m5BNcvXgkFVTBFJJcUtNwucuGvv6cpjQ7U5tRCMk8z9iGizAlKHAYKeUT5
DI7h6pD+GNfIzdvUL9w6LuMiI2zjuNIClXCT6AshFO0bXfManOpgQk0/I0QlOfBcInKFY3oSzwmX
7lNXh9aLXOmiaIh51F+Pxj+D3dLeaSYJ7Dk6nW69fcK5gMqNqeu/oT11ZMTLzZmqHvOOoyWgQE+G
6ZmD8EayNzmGjL69HVoSSIU6xM+PZu+jkURT22Jb+YhroRqelxB73nj1DMu6A4D5Y3wXDDvDwlQI
XOpTQRbyCkSgtegH23wZzt+XdtAzrQiS2wY44tGKFfZtrW44XFaLJaIlApeVnvwhVXodOJ71Jrjf
A5Zr6lX3Y1CP/C5l3m6x2atCZMZOM6Go9iGcfvSZyoBveWWCAuHGyihMqC5FxGWQbHyj98/sdBAs
e1Smd3HA/kzezDiZnK1zXCrOZI0yxFcfgS+ttul04tDvoAB/2ZO7+fZYugq1Cy6nOgmbthFpy6QO
BLFFPPHIVPe8eO+Ks5zrW+/7B85OT4trsZo46bdApORQm31Rr5YVyuPIHhsQQLWCa2AXPmtRhOwC
UeKPVlmjc/s+t9ZMFR6ebH0FGBSp5GHIOeGRq1Vcq9Ly70uuPjvplkNI8yJ3V30wpqh08yo4AHbP
RDdvUuwJCPBlYAo2kitmlvX9YTaquzMcqMYozJvn7WI2n2mqAXvHuY3IOSiPP81+xsrwSAqAVxsb
COvZiII5EjOC155aBj3xHuPR2Vc8T3c7ECOJ4VGlQ6RqFnvO0OOhR9OXL2nPH1s8x6l50IK7Luhc
Bdjzkd+CCOAZcz3eqHDwB2xVITluSZIcPYtFsK55Uc8n+H/U0igPU0ukJTq9qAGhcS6zTa4UnlzP
Tfgknum8JSVHKXDxJe1V2KbdXwaUB1YyiUjbv0DrTuwG8ddfpWZa0GeM2IARTVDk47fQrpUO7T2w
7x170ctkLCJEcixygjXhTPq9Vg+edaCanoo8U4J1y7oE3C0p9HOLn38doztQKIWd4d0/6XW/EOPX
a/kOPiUHMLJ/VX93bUWu/r5oUUtOj6j61eP/dzDDoY1/4SgeQzolyNbbVI7RWiR3c5uRoUCu4pbZ
ZQSzvL1vwNDs/MN7NK2iVGCUfDVBK8gEa3E8gtABmQhXMYYnrWDGqJIyEV6UfSG9mOYKwH8GRacy
WP0AxcZM4Caog2cn0BbqP77Bb9B/djs877oHln01xVL8FOkR31utdd+8sua6Ys3QGa7mfhCweyGM
t2vKk13e8uawFT5IqLJ0AcmFyLgKPsVibXNYbeBioYVfuIojod561KXIBMCeYypdbO/OxJ0pL0tI
c6M2aEad2apylx06ALmI9kqsGXo32xnI8zGaok38B+t1q/HkNk1utPaGZj6TH+bg25be027HVzxE
4ewj9nwotdpkqsUUldYFgr5OlWSlfWK2qqEei3qsyecWmUGEVPROf4Mt5Jo3BB7xrsZ4w2ZMP26f
qGJoQ0cxgBKJJV/GyfM6UPb+q6dP8n3gw72oOx5+HGJIHdagBAkMA4uP7N4ckm2EHWrdlkwsd4WS
7PZOVWsQSNHG9K5yBnU5I7WTRFFcK3T9OByg6bTgrAubYDYqmI+VwAWPLfIxGY623oCRdpi3GV15
nr5rfk0z+5KZIfZwuNTnGWErnnIJXjp95jOyQ2sAcoJWkGYht/MYWkgu6nv40vZAHPqcrjm/3g3t
WE4tVKot1g8x0BX7mpPU7njgWEv26IkA7jK+eBs72iNIQFPqJ+2kGX5rFj64Kt/kQXSV1xy1MJXQ
fS4Tdow2PAVMFqsV/Ce1temojETtiro39HbryWx16vJg+pU31jV4p1yapYynfQgpUhuf8YGWit8r
N2KWxnAUskndPRVCrYLRH7LXR9SCEX8KRlCfS9+7qvJ4AtC/V4eunIErg9NHUChb+Y0lpx073e7n
FGKFLT7tfyaH2lxMaotrMbIZbQgKiYw2aOBvb9eiWhCUzRenI7gpcquVFZBJMxxS08FpJEZH8jti
YRYcz0flKELj7PSgu+yfI926g7nGty8wfinx75wQaAUj6reT6JPGfU0YhAfBPJ/8enkK5E50gfrk
qIZ+ooiWjZpCh9yXuZPn5JqO73YCrV5Pepe5sBJEN42mtIhMYCNe1vH65O9P3uOydfBVz21oOhyQ
hBM7Lsj/Nxyb51Q7uvvVJzT2i5EfZnGzDWXYuo8KHC2vuFFU7suAZ+UlgxDJ6BBoRpjkDCuNkmgV
Po42/kA6/++FnAr7Mlce9sydEJKy+TM4+E7zqDBCC3P8Yw9dtnfYhKKjt17aJht27Yz/Fen/5jW5
UXqBMtl9uMEejFfFqgD4soVx3XKtRc99pKblDtbkrft1upJPqeXOzjHGRYqYvb4r4mltyYmH7R/3
yIoOGT2NZTKoP54xJtBnlgKVfz88fjtzI+eSIXp8dWM/ZgkpHIraFV8Efzmg6TPGDFS78apkcnDX
ML/p+B3vpYE0I4/6xstf2O8uBrjQAR7Sw8CJ864iiJSeN7ab9pnJU690ft0dSH/ToYE/q6Hn2IPg
cx3J4QnoL+Bm8j96AbEYMZg1knlsAOsplj8iQqv/K+bpZL13JkMcqJ+44LUAUcfKJmNyw5lJbjwN
GoyRLPBJxuvwJ34X8X/9hWO4jsU2CGRnrzM180gDCidHvPhc1WVoYsXfLOQPilbyA3S4hJ60jWD3
Al+Na+uuWKd41qDksiH3ysFWAn0aELFkOsywTD3AjvMDwn3rPJCpf4w5wiuUhAYXV3Nt2n93ukzh
TdhcrF5i4ZNc6UdLH4lwKERxGvDCjhTLwmzHMwtyrMwDwyVd5hbOUIho7uxfxrh+mezBBXcZvqeK
5Ak0RuBQOmpIAUgBjDC7eRUtURLR2QBlhYHqFKZhXTFYVYiCVmIiltmw0NbJ0tT0hFF3R7g99zEH
pGfy69rDKx5YajJyrqjulGrP4M85s0FE4oATPQRZ4wxTeYp+XlYt0UasloBMJY9++SEkkxb54w/c
h98afoDQLBL7OgCzLVTgI8QIJ8Gpz/8AWpE8OvOrdfloWUH7uyXmw21NS5c5TamI39hQvgWw3py/
h7B1cafqQZgGgqB23NfjbgooAWM/3R1E/WStKhhecs6BeI3uzgczgF8qN+7/i0iPkLOE8ZOTRljP
5qJDBVqaXWYlqbJ/h4sspEIu3RrAN+JgzsE3ZrHEDH+eb3EQRpMdV1SYCjO4FIcrN3hSLR4HhOUq
L+DwHOAAqP5QX+225Py4cN0UXYATX33XUkUqAG5m5aaVInYgy6fsMo+HY85CwRCo+as+MWVesQpu
jNqMIukFzxFq/IlBrzcLV5b5975u9wsj3676DTGpqi00bMsDm/gDgLzLYD9Or6NQdm82+ztk81Td
1SZyLS3t1DWtCn9sifOCvjpA8C3W4hS/57xowzMp0vjdlTZGwjTnbsV3eC0fu0YTNI+gEYsiZR0Y
nhIPrO60Kd5h/jnagn/dGszkwZ0UqLDGGGR4fTAaYv4CeuTnSiEuXzBlzw1/Jo+vPzHHZL5ZoeSV
ilx2v1lZfP5o3E4RYui0YOFFV/C6WC08ePRfxw8nQvvKwOnwytip/UO6bWu6QoONBfygg6NjS9HX
e7Wd25lturQXqEYEaJ5kcbHaWEl3J2Wlf+6ZgDjbu5NqEy1yD9p0V+lPqwXyqq9rC6rmczCsqNtt
usMunefMj2zzQWdzDaUlXFdHx8N3fXEWw2a93kbHrn27Ga7mGtiNoE9zn5GNYo0L2POVu3VcTOnG
qvsU17a1WW54gM2On1n5q5vYGGNvzCFAubd3SeadGIZeGytJSDOpeFjwzo4hHfIKuR+g96NYOvRR
mdk+DI2DktURPCr074X3XU++wvgMR/ZVuFEo0hhK9Ea8NFq4BRcVQpUP2rhR8XlWtZ+Bg16ssvcz
1oX0dAIivY8UtuwcKcw7KOUPKIExfLbAD7jR0k+0yYFrRyRGUTyvNt3HqgGUl9g/voByTQlcfo2F
aWWTgBkJSBVoSlQwFiMwVzD4nZ6AiT8UePNIQtMNmz4TQCzzip7Jibxs4kGq9jOmooDVerBLa+eS
q5PTOTSiampNtemcs5i7kd+cTGkTpaBe4hUIU2K9jxjpA9Nx//QdMwhzfCyYzS0BtFMz89DfvY75
wCuwscsYGrBXWlAtCvipeBQ+wQPQsTGObQZ80KzUPxD8nGYXLlfSmu9Oknbvt0NuOmUGFSDLOlFK
V/eZU9wNV4jHxNqvRyKwR7IJT+IIv9R6LxzerpGDewe+m/jZ+LAzUXpHcLMCcslyj6aCtL89nklF
wmEh9g5Gp1cTcxbeLMExgvNUI+vv75I05IJ7jibp0isRHVbNszdn3fSg4RyfpC2eN/Cg3Eea2UlH
vMmYviCbVSweERkWdC9WCxdKSXaDYCAdUqr17HQmE9pFNtRIq/IZiV5LunFMTWHp7ELcm1PSKEZk
8/OJzrDox0WzQuGZWtmy7n31P6O1g55OG42yYjuSKpopIghwcqwlLY175UeVHY4u3rE7hDGfpJoN
UkJ1+xYyo3IBUciydYjMQcemoAcXT8Ol61zgPWDaoOElm9BCiRq7tXmk4IuwJQgUKZkWXp+YAOu8
o0NWuML9ftAZ523kea5dt/UnR2kbfIe1+CI71gjdsisM3489YNAa8lHJJBMASQIqgP52mvq4dR3H
2w6lsQjDVXRFSgWCYOqip9XVgjbroQNAEhRy0AvpTqG8/9YstbDBx2aCUJmmxNYkCDMXJOTMShzD
weNuN5mBBjaXrRMQIi1zsBUb3CL00hvBMCP8wwmqKTLdDiMSz9KrcW2CKbvCFzWRYwm4o9LV63wp
0rXT5lGw1TbnjmzYxdoO6pNEPdiQ4yyOY5tQ+ROBqrqwhIJZAoMHStrHnsju6bxG/bWHJaZEMLtT
6PmNvXkf278kOy/xPNaTxV3A9WKoXAi7ybKu1xPHXP2UGgi8stjE5J5rA7enHxKMoTzaJjr1T58/
u0E45LRvCRha/EGK/d4CJDE4dB8g7yQwUQGC/se5e9sOwBgfdWd9eCnfc7RaOfkVvCDQAgDZdKGF
OGFldBLyw5wE1EZUah1vkPm7xsIZvwOwl1kwcDeFeYUKkaf/+j5DHpYTD7stdZnUp95d4zxsfS4R
tFREzyBv/GtNvECdN2j83czIaN4b+f/Xm5fvwVoFneWumkcnw1ex65ZXPWZpM6MRSqJRSOKQhWjK
fNFG+6DUpwPDGMubm3TJD1oniQjo/PCzpyWa3yaug7I0MRTQsaPPNrWBA2qEkmErvLvlOuZ/ebm0
bFFWiqn5U4ExCldl+dZp3RK215NTwfTeQwfFBPmd/uCIylSrbpZuAlneHL0CPA/EoLpeuYJ3CM8p
Vzal8FVMqtYETqrWPLXHQXGiZBda9aCPaIRP1+LBKsViGqR2NtoT6Fn6LGVdG9NJXImlcZnM1W3q
tHYdiEQGygOFu3FrcCcyOn/kufmVdQ0ZGV/F5XciT5MMYw+zedlyHc3Xe8GJAmY5p55Fw1jwIdvO
i6gjAGdTy/N4/jePSdGQI+nNLlVtCD4iif7kKcC3a1Jmfr9AynWQcbgvtMtNrQXQghY/PWAK0wQg
ujLzTI3FDq58YSq9LF+vLG5nDaEpwOO2LHSXaLAyCC7HRXafRiQhobcih9Xd3lMVLdg/fXCE8BVH
aktusLE8XqN+W94rx512cjFEjFnGDMyizdJO4RXsu7JuZ1+gDkeeOEk2IzZ8i+5NRkRDxit9RkDR
cgDh4quuPEq3Oo7mgXvWFXZ5rvOpJ6ScqyN3riJRWc8rQYJxTjvmo3u79eglRPCA0Fo1z9M65VUN
6fPLgoR82SXGhgG6+8SZkMwkGF29SVVY2xjY8RvU8QvIVnvxTJ9Va1BgH9HY2Jd5ZZaPJidy7vtp
D2gkq7DnsjYbHoUgcaUDkBE/Mn66/qBW82gH85rMfiN0iwbEQj2EPWn/UAYIpJ6kl3lHqTVau48c
dqq59nR/rsT3KYqO3c1KUzKG8eMezkwZxq2CHqs/Nkyfrcnfxb0lJLJKVUfF0Xf9nTEjcRhKXfGQ
2v6myOEzjc5YACslsZWg8Yp2jhazwovq4kYNO9gyGXm51Vlpx5AysEZ7tbdmSHA5Q2J3jj/DSY8m
GBU+4gLqSM+jwotiP/6+LeQ9qA4pZuqyY+zyX9SU49BHpx5x+sKVyXvV8i2co0jdeUSjRZW7Bi7E
njP/N0G5kGcnGFlYb6VQwgyl74JXi6DSn4sID/KGO/z3eZzZDyOGKNz0rewelqhA95CSCuNH55iQ
vrtq+FVOVQMfocyAKAUAsbdssQiviUjiRd5Sg9KmA3uslM+ORPUGVaLPkgKZ1aysCyW/fEu4WMcJ
D511qSxGfqthuXDARsNk0/S5B1sdkw8S3oSPGfB13dc/NVeKp6d/dT3SqalrTjODhiri1cC/+xMW
XwA6xBYzfmXsTUe2dsmI8EL/qoimaYuEdaoYhKDSVjnRabtQsgEhb7Tbdk5OkO+moPfzlAOupOTc
bki9CDvq6QiHCe+CmQ7QwPMMKmlkBuRQAKd8s8S/w968nChOhB9IHEfhYojMhYAwO+UCBH/kvqAC
jAkqrkg6mVwaVBLulBwRAGPmH1phcVL+AFeVeRnLMUhIeOhKKSmOAOygl3LPNZJphC9HrVI7ZJcP
uhCoSG/lX93Eu3wM/cBodT9ISXL/S+zxqxJ7MCR/c8WRTlBZaji4tHHGXwbNiJvBmC9mIeMVaoPs
NalDw58lflLdREFdHodUYV6pKyvGOU/uo27K2QK8w3zs/VLoDo7CMFXLOp30TMF1UrSfmaqzh7ta
fBc1Ze/d2X12OuJCedLNEaasqI8LRio9vXPbVCjoz7auvkLbJWBhIm2Q4X9tZ2AgFlo8OVj5TibV
VpcajE0ihAQ3ZDOhD6b9dmIGSEk1IITfZx5CWRjWq7DXtvWbGeXxFtZcXzqo2S4eOjFdunMol19N
jkjamLvjCxOMb2/iQk+P67POms3p2IpVLIx4yPejCY7VdVVPnwNr4HZgJWrMSfppyff4STZQyzs0
bt7jg+XJ1j2aPDHZNPWUtuJ9dT9csdZNvAlBBofiytzZw+M3b8HQ2nphMWNViigQnq0o6Pnee1uR
jnwaZuyW6uNBRQtkP5kMkm6Ebl9KXeY09d68oFmM3azk73aWdl6R6mFoOnuTRj6VuAG4Sj2FBcQT
wgArYC7suFNUNFHCkS50jFK6hf66v2Okjxe56R9b0GffkvdCJuWCtd1xc8MCbTG6RoGm56rQoH45
HiWpP0fEi7C/4YFrykqkkqmZEhybiyroqKrOsFp/izVWTuWCUNgHBxGq8m+bCgh5q+FTk4RoHXyL
H1UxWkO3fs02xKZdOlyQpE1pNbNIQN46OFFojWRqi23d5oHQAyY4dMZ3vseKR6wLJitjcp5V60VD
15CYnwhL7rX/ZFpGGGS6CibgHDvt61XCEGuE211VE8IVNALe6re5m5roAmb8wOUemNyHllcGg8W/
xEJXxw1Dm0ntE8ESBXZXGnkxmaEUi4nngzUZpUwMV0YP5b9DEF0ZtUoKI2znSgEZQfOoStUDkU+/
QTFzZZ6w07BVOezmIuXSZrs6WYWV5cY8ZXnwh98tvc1iqYmP61prwY0M9a/cspYp8WNlvib7n7A0
FBSU7HWm8oVOt5B8CO9G4Yk4+/vItcdrJiPo8oowEBuudN3Whb3hBZ0RNtlvDlJZEg0YmhK1A/Zb
qJDek/hKY08YN2Igdz4QmwEcwhePw6hQeDADerwtE4qYQvtv6yxi3x54NRkhZHRPXSNPOyUSp7Ij
tXn0ltaJYdCEPC1pNsEItKjbhPd311ObNqxOeLFMyhRJ/UVldH56tIuviZtdFUJ+fLpabQHjuBNr
ZmhEe6+jL/mkR0S1v5yHquuTxAiel22244mif1jaROVyWLiyNRcRpi0sECNBwuuUIYt52s58vPdi
AJNd0WjMw88Vgtb5rltaUh2IxNbOM306ZLk2CscNdW8JZ49xf9pY7uDJ0AI9i+H24tvjKomSIVqt
mSM2qQzNKpZMncshItO0fJ50bfIKSuLAQaREg4pJEWNPB5wYohJKpCxUcc+uZwjTwZdzn06h6OxH
Y2diA4z6UrPsvrmnT6OSyM1xGKk/zUAvnRC7dvNuTEOyD8yTYRNOO8Cu0ZdTsehrb1NZQKe3mahh
4UBqr/5f88skxgu2jiQXqNCvHuY1rBuDusB9TwjkICzn51awMOkzhU3xrJcVyrsKpQtqBvuE5KD1
+y9QHkWQum8HQxNWlHoaXxkRj/0r4a7nBIoJ/Z+Z2T69z59sQz7Sok/ftduZBWWXvnO+GjR913og
bfirCB/VOsno22rHtQTLEbGKH+eE6CCrV+cFdLj+mFU1mO+AIh8ntVEWzZQ5qfHRTCYZbjyXo3y+
ygBo/7CFN6unxiJipAaWcqJzWJD0JMh/cG4RGDFLLIJXOslRjg4Ep6vts+Y59QtuniSfOTIrsG3P
MZ7+/EpeW7y5c5icoKVfBisyU9mywxDR9x1ZcIGp42X+ZN1aVr6BPEXnzNKIqKP8os5jqwPYXLHV
CUzcMjsdyScycXMpGYJ7LXzjqfxZjL95lZbn0T9Q0KeP07TOAI/Nk4ej2gM+Wxvj3K3opHCaC5nc
7xREtK/CMtuqFXthetsPyYaJOD617GgaTkN/tRqLxlI/TDLR8wqnfRp1J/ULHZShJoFcItFjQ15d
bFIaoZA8Yi07h8JI0PQTbafyLXKDHKwgzM0WOLCBjQh/kwJEIaTYjzN6fSM9u+YVhxnW2BB/bCs+
ueotjBaK3I69/Lmd8JIRGbcaRbjs4Xa80P7MwikjsbwepN6gUdBJUYi06lKG2EnLzlxNRDHmdAnm
Naz3oNin00BJebCdi7mSzyll9zx3QCK5+6vK82I0Q2zLvE9Z1+btYHHpWyDM17D9QZDVzHL4TDwu
6L/1EmlRwpWbI+c7QmyZqLu8dAS3l0c3m0XRHZKM6YGtrYiBJaZ+8dlAiWUqyDc8+l7kYI1XtEyI
jVVOxon0p3AyJytBRaCuFY6xpz0KI2dgr5szVju31v1rA2FhvSijvi+f3HHLsAL/dE826jiQImGM
se0LlLo2bv8AmsByaNkZuWATQHhYMpWmEeGfVOXn42dX/h7fJpI43BDi+aWvrOPuuy+/Z7+ctoqr
pzNw+kZDg+UvOSeP2ro7FxsxodlH+2HOCRFR3DdLVXb1gOedQGzwsoZBf3nb/Ub7P4S5UUM1Rf0o
me4vJoUbrpmoVBLE4P7AXwaaZ01WwXhMrxJBY0vjxnUGdMlF03hnsibV3Rr4dibGnq4Zq+ibb5pL
rBBdfLizkIkhn3tqsLMINGy/48qU86/UzGyvyCWZu9xX30crXcUn+Rh4bkNYyDLS8JgsSmLMUIgo
WvCZILgIJWqG6TGBLienu5ZXLMuDYB6yaG1y5dcUzoKWfaKQmXmNGpQnlmC0+fn7REUh77NFISbV
wHRX47rgq6BDvH8cmPBCVPTNJyV3hrCycrqwJjko4NExMhv3hjB1n5CdywwzBGZxrGfEGrrPCq+B
/HV4PQ0OoqgiHnGTXKoxW4UJzhFgyd9rQB4dEVx9YMJwCHBtFPnV1/op/MPvo1PkpJ6dR4YU+EOp
qE8i6HiIil8yMtgXqItr5f7t7BLI35+D7g4b4cut+WmbSp+nL3t61M7XRLFHiuE8dnRKhOdfgIRX
p4wYIkzEenSbtlICalwNU/8LwkgSG00B2UO7gWQspLHZ9JcCGomqz/dvK1wzuz7PfmZ6f98dt36J
wWh+PGYRr0TXBI9TgX8ZAj0vZ50lzXZgyL3QCTeHc/b9if4C0Qmk/ggT4DnxVYXm/aBtyB+59GNF
M7D58FkQA4bFEkFteQsSHMdQJTVVxxUb+xG37/iW2n4SoIXlHI/xUpzjZ/zUTZoBPa7tRH4cTGmc
FVqfbvu49spnY23UH8uSF/cv7BWWIj0u1QnP7VgaClHFA0MHqUV39yEnFzeYapMpVy/3yUnsklxQ
PADbgkNJYfKpkjMtfLbAWokXKs40o/1TJITuQMYEimehdGfw9+13GPk27YlY3l+jD69cS8HC1prn
L8PUeAFxnRScdwiYKqSrV1vmRXKoZ/WSzziBY0pq9CrshnhEb6b23JIA5GWR6dIE6j6WXUbH8Ui+
sVpqDTcB5Qd7UKauoED7UcnhpCeHsoBKVtRCI47mNZ1OAq/FGoMfyinXiOwPirtVY2qZF5QEWQcB
l7wsG4eg/PUzHxEA57Ric5aq2PjFsLG0FXChAZC/gCQ5wRjR1d2X11g5/mKStZhqwzkyRpmwZgFR
oZcgcqYxhYnX7zzuVL3YeOG9Y027DcPCkOglP2PKDr98jsPzj5+9U0jmm29uTNJyn2vty1z3JByw
Csn2/E/B8bJZKj10j/nmo/lj2tIFX60HQ9XDVGOdLlRD+CGGZJsepGIdgJyItK/vHSy1kmhoJdL0
7GFwUVvHmvNjcyK+NGXr7yeevzg4LzdgDgyVtU/BnBJfEAh26vQe98D+v1Ey7B2NkPyp4Px8BxCn
vn5sEwVA3GADCNhpuSicSgOtqffNGv+OEwEddsAXO5Ys0a7qGjRos/bLk5aHzlEwZNYIIitHz+hf
hK7QH13YRpx6v1uiDpP49Qy7NM6bFcH4u/92ofNoTnr4wGU9xHceeFBbufvx2tJLptCzSUE8dJPP
V6wUJ4IdRtYWykcpAc/X1WvMr4j8a+knXRXX/hkZcKrx1HPOKaz0xk3B4S8JLdZjIQtjHk1mE+1y
JykGASQaNEd+75seaH1QjjqKJwDxVsYb3smbCkEBt//rcvqTlybYsa3YGoQ3PuL7tRBbtMsLPV0m
/y0n5iOQKpFo+X67cmQX9LfiYhBsjFezbth3EC3EQEZHfI06kGKtlxNU2kCcv2CmsGwtg/IRFPQy
EDRZns2MM8h3S69mQv4jLtXaJpKTs0GY6vjbVNOi2YS/uvcIeHEhA5CEnrduhdJxBL+4Aaa1qoRa
Cb++q8+Id7MCq2ieD9ACOtpMnQhpwvCOmgl+VEDEekqw2UBaS+hJG8HfHEMv5oKzncnh4/B3JgMN
0CgLKEQa5+23ydx24hss2Jya9jVqSxyDUtm0dGveovcdmh58B/4hqREBOt9WvigNAKRl1Q5Adaqf
N9EpGlmJs68zYBxtwa9WSWy+W85+iAUO0QUushQTfUmj0YRb3MmwKrPSsCraxcdu/xCulkJqYcYg
WtZNsQ90D/JSVH8/sJZ88B9/rs0tBA2/0kFnu65Usw2XnMIN/OwYzwWRblDK1MR5ezh7mcM1Mxt4
H5ujC79eXJqNiyspEtesNchy9Dd8vGkMiz40Xunj7j78zMGy5zZJV/twmrguBtJXJ7pTWuZQfRk+
xkQ4FjHC00lJmKBEpR/ORVJxHiEf2S9zbADGnuWSYNzFc1gIqDIok5Hmgcc9gZ/tv3Vduo2i15DO
ALQuwwCCEQLV+iBkPSKy4B048mevvGFAIp8y5Lf6kPSNmthn4rrL1q5BGJS4kTqLMzo6Qz29lTnz
9a1CE9zQlcFZLdjT4KguuE04ciEo28qQSHscv3C7uMOlTG7cTNs0yOoVUo3LnWSpzHcvIuxe5pLm
6emNRNj4UCOw/VwwE5VD0c6JDUivF5PRRDl0/O9TH9yY8owS+5Bf0yCtGi7dFY21yII5gB9TsI9U
FVuFh0mdfJKirP01KNq53ZNfAI5EIi+29SBEmH5y5DItDcIZeDZXpm5E3ldSoyGeApABYEXvDIpV
P++/o2R7xGsYX9XVAogK6qjjffk1haFY9S9KWIK+qVmlujHHJPyXqNAZo+MmqfJzssdVa2URCYNc
/mDxyvjN9XaVBw8YY9s+VK/nlqUocKdDsnKPhYesdYu96H8oDjMjl/XWGOtfsRtlItM4iCaAi9sD
Rwcp37+4AN8J7kKpImKDHmhQw2n86xMl5aIXkct7N8cLbNwBofQBGfaYXIzQcNDdzNZXoigzE1Wd
A6PhaLMsYE0bUoamFLAnglYRnTtF4S3DO+Hm5C3QrLzhQB1BpgkfCtHd2OBLRa3pUVkGO1ZA0gvB
OfHYs/n5lzu6Ox/GtBfQOH6KnJYpS8PnVrVjb5FlXKplMsGGH0Mb4kkRDMpiXLQ9bkszUr0bVLpB
BnaaXReQzCaJOeyhm/GlImi5mahGAWRgEPxxHFqeNdWT1Wm4W0gT3yPuAN1alGHS6BxEye/oWw95
PQDqeew/J2PvrEqGR3oK3f103BhKc2bHMwGdQedDhKxdaNDGrmKlLROrs15RsKRNscivtigx9kuC
iVa8mN057Eeo6qZTbOxxPt5BkklirwGRGtFt1anjy8gUx/RpKhT7ann3RN8CUMYIZTlCiqUzp3MZ
avG7VSUO54aJxDE6FRvsdvzAbaKxIkM0o40gxreBKs/gsxFxPpx21G2NBrgjQ0ck2wJXHwcP3iIY
i3NuP/R5xQ6Pi4xrEIYceBrhcZKqEDq+SOTo9R4/9mLdc421DfMwyYMAL5DQx8r7774/DJCjd2Xd
IFzXE2UyUG7n9aQHcVlHcZS3TZnoYPsgyRxi0AbReCF1EAKjFw6rjFBIZWBDZGiVadBrM28MjVbY
znzr7crjHDTeiFTE4VXu4JhOLKH8Tt+xZZvtYJiP6VRsriRzJkFzjNhf6f5YmK4g9X1MRtgMH+eS
YY2quq6cnfFUWjXiRxe+1Pk1d9TXtgDdt/sRTbHT7H8TIYbc3WYQhdmFDx6U3FkrUuUl37ix08aK
F0CI+9Rt/KErjObZ5U2pUq4r4ClxDWtkUK9PIMxkjlDb24/WboLgq6kTYkdnfj9s75GbnHEQZCYX
/w0Le0cUoUSWNN/0Cr4pl2+k/veEbiN8WuHLLS/L4sKCIkx3jpK62JULhOloNSKkeAp6n9uKRyHH
RDUECEy6f/nghPLTysuoN/iqUOQQGuPlsvgTwqsb7VZ4tGvrDHXjjz/Q+7BhfrxwuNEwCeecS77r
hnRDqtfdTfKlz+L3va1ip2LGiUmsxnqMpfPj97fd7f6TjKR4Plmo3Z8hKSIdqC9PsIagvwkf4nnM
slQlxHZ+/ZJ4GD5Us9PdwFmxtbjYL2YrgieornPnTSrgZGOV/6LeN+2AkYZHP7x0sMPTOnvQA8Of
t1bO9gWDRXHilpaGGq8ar8RLzme82fF/iqEUdfpqtNXBzN9R5sQ2zQOCysaO/ET/PqE7i6n2TVOe
QL5wg7RUPJ/4vc/6QPnAXhahNjsgO/rHq6ghs7gcx7MxUUUIy4yr5QtgXgH5ViVeGXSCDG1LSiGy
LXMuGliiwmRFOQD3FvFylGPlhVdIfkVcoAxZnig/5DTbyZApZYs7nPs3N6MBva0Xr4shNVBYXrKj
0GIFfS6sFYYftkaJYJyNBa2AFpxSMcgIVhXMKjPsuiCavWTiOi+2e5xgzEFDzVqUAPGNM3v8JPVZ
Tm8DffghPsHubG2ptILPJ60DY78evkQ9G/IXGtHEHDvzbxtntvc+dBtZAlQqnX5oLX2Outg82BKg
BUDQx6eiVr2sryg5B3qd1o4epR+Df8bZXtW25llfwoJFFxJc3U/Mlz1eGKqT60Fy3FDAWI8WtpDC
Qd2dkMYA4KHXQSgHGBcDUCl46wrA8l95DDUx8r/Yg1L+IvIGxlPsQqyziEY8azjGCEMI9Sl4nNge
1FyGazSBaphRv6RdG7r5g8MEi021+vNpIM+b2CDO2TrzVygTtnge4Gz6HFvXEZ1k1HqHmS+XwL6z
2Z6zbgMT4VO4CZRc0Co8kqZ6uDLc6yHxXRIz98DQNs0WLxpogSKXtqw3MFrIyv2XamxITLIFs7Lt
ShLFoetSCGSMCQ5cYOm7eb5xzI5cAbG7D0vmJkBBJtfVjracWNm/1jA4Qtq4OG4ALMpXAxZPl/Qq
0ODamHS5OoplxejlmpGBpH8zwtJfbotXDGci0oxvaSjjrg99J8AF7I/qpke3bsTwJqAxtgsU6GNP
/NnA81BqcJYtqVXUDFeIcypVXOyaedKdhjMkTF6LJnSUDlIlM/zGstUHfNpPoX2YRP2ibxgxDkkV
yLkTjFrGeoVryO5YdDvtaeoh/pps1DQ7haG+AFhgU0KzCwjKV+kcoiNs8DyoB3k91APvRKBQksDV
IZiOPlwyp6Ov0Jzcc66rShVgkHqIg25e4Pfpbz4dKHE6eOjA8nqF3PSSePqgufsFoDQMfSltJ/FL
QaxLvDcuE5kqrnCPdmVSRZqacAejpaDoy1X2KWzsPuwA12XyLGsb+UMJvZIrkYzNHHgWxpYCwnFM
bLz3m0Bs1998krJHN1+wlXkZ0xr7ZQvmCZaI3WV/Ekk2SBk0sMYsc1BjzQmr+BDdZTQ9Vmz/MMa5
JH2dAZPsgUJyWrGHK6Oi0YRRl0n6xJ89PouUCRPcKJ3j+/dktlZA64wFJJQsNXnOtLfpEj6jJNHM
lBIEn9eRE1iBiq2RvSZpSPtPMhmyRupcPUUz0wuYuQEV+Useyn1k8ZpejjAK4wd8qirwF3mgJxbJ
MvX6KoEpnXSIxSpP+4u6t//iiBke8z+wG4rAyDP55NVXuWlePLYSF/DGimS8qx5gTnL1tJgjnzoy
nwFxSXYMqWTiCILZ9dqQKQjfplHL0WDl6GcR6rZ3FLdCXyrL+Pq4YBhmX6LcG1DhDz6FpeIojWqD
D3Hp038cmkrigfn9ZaODTY+De8hmirqDVHXY+RWb8Z0OfM7mdiv1o7z5J9mzru57wJ9CdmtjSIos
IQwML+vv6RzyvdOEnkdp+iW3e9swAEA2/UpqZ6kC+lRzQNmhie+qndFz4sGpv5bB6Pk2x/VB+Q+7
j1qNFCvArJSnXIhxoFfHbXt04GwcKRHau84VdF7iXBmEp+FtmXK+TYdFXiPOEjIERzWh7bgSFUj/
nVqtHjdjclapZUEkMmPfDWb1B4yRX6PMBMsO6oY0Z4ZDv3B9Wy/K9ypIqANGAVXwKtOZFEwEeR9a
H4u54CjWz00FTek4FHba17rX4wvqRnVfRjnUQR+ifTcYGorXNzsJyzmX/XUBnH+uzyzpYbHhLXhX
2V+O/pGDlKMmW4hFn8pFp79EP5Vng2uKKUTJDkSCMmDpsPrj4FQ238P1F4m/BpXk0RisDh5ivcgY
oynuGuMdSA8fAHdO3bJENonRqYGTisbO9n+htnM/YUsE3HuAL1zSVJOLZsV4Fi+WcZ223RFi4WQX
4/Uz2tHBmOUBvLthYhLkVi4shMHe8IxZgb/kItTzp8aSN13clQp8k0/sTlreyA2yYCcAGHCOjvgB
ecTh911owZm8+5DLHd8FMOW3Bhuvp2q4xJIEHpfKi4TqAXvFLuppjQgccKgwV0WV7VKGdDYNxcaU
vgbtp4Tu4VkMILX/NKUJVF5OMD7IvQHsDrOaO0Bv18ouc4spRjKrdRccZpY6n+349OcGZ5VGUO+a
EPlX2/HO9gaPwpAGl4x2NY3Qn0cQM/2v+dHbd88a7uQGsDNxtBNp3pkUMrNtLZuNXrEiUCTzFS07
yy5xwM6JCLNihKX42NLXomvB+E4MGcPSDcZtK38HRjep3agY6D/ahASzrgTRZYTbYWd/6H0ouUes
09bYatnA/imb5Bon89tI97+WUrLWmBjQkvvpEAOXdPVfF/EtpA0qC3OYLc7ZmVPLl1UTTnEGyR8z
rDv3/6FIVbmgAUukA0qIIe5JJAnjS+StTG52u2AqFlPa3hc2nR13K6bKepxTveX/W6VDaIvQ1ISx
D18o3jcK+9jTNWGaLCKghfbElw+prZIAMbgmVoj1G6IWuu6ecKw3uF79HFkR4PWdapqUZyvfsunh
ZIePfOQH15RMi0qpejv7sryzeObSaR995w0/p8NAUyWlnIqZDDg7UZke+wZqqUF+5ytW4pUPD7vC
Lo8RUZFvc/HIr8FksqWqosMZnQSNNOjRJUEf+XQ4Iqy7JRCtyuITZ2fvIsLFPem+BcDhigZOw0J4
PjmKSMvfSUFv9RkNMnxzVuJjSPIShZ41oPag9vnjtfuRZaeSh2wRi8o+QEh6K2VxtB8obXeGq2Jv
k1H1UJjvPvZWsH0eI5P5imQVNt/rxA3h+PdiG+W1h6s4e8cLoMftci0qdJXBnIFyTecuGp1QMwLf
+78s2es3MevY6WPtnwWmSbbTpecYlQeBqbjVN2+ET1MPzLlC2/MmJaMJ0vBeOofa3WHUpu/gZ0bE
WcK6/srx5c7X/M2NkY7Rv+S052b2edI2gvgCbYjBVTJ1w3bDflmGsw2kffweauol+hvCAhPpX8se
LdiHEHJDADYthUnulmOwv9YmIQTSPCEB7TXhyqag8dufT3zsyAFVBKby0FnUYhlXiRoxz5Y77iPP
QgowhjZ9v/8W+z8mTw2yE7vRKVa4bVFHtkFpD3Oozv98/GHHXqMrcNhtDGuWb6OSpmJGzc+F6lQ2
TBgamNBk4QfEU081ppdsYoUp2EH8qqaiyf8mQLvezz6jSTC13K/GYP7pDoI+8m3Hfjlt3zbaJoqQ
dNwbdRSLNMxRI1emoWIfNA4TlSK8RqT1D9327U4i7HBIXpgts9ZiLiPrQLavUbzuY0vSEJq/EhuP
97f8SG0gLv3uONaPw1HfYr+1DvLk8YqmUAhk8YzYYz/t32b6t1x8EjXg1G4IEMTF76NULCsNYSSZ
To0qCdTJR7VFZjYU66UoBgfIFKcsB/UANdH70czFnUoN38V36Xvo8FmUeIcXAnpNiyt5kYHoYv5/
gPrPt6cuQ0rQWx0cRHDxiWzODetJs77VMGiCSAgB0ZXgvDilMwD4yyWGcdj4wlMuc27hCdXEWzUz
17MiVkP2opEQORje4/q1mxbRHbuGJxCTZT9BHIYJ16ODK4wATDIM2CkbYA14eHpCInORY7MyiTeR
75a57jE1l63WKJjxyQMBGucclVtQVJs8FlSAhFM6Jl0a6Qjd+D7VZL9NMFekY5OHDV5C4YqpyStV
IiXTeMAahx939+UDr7y5xp2cy6MkG7+/MLI4uVVfZtqasxQwFIdSu1K7Wt+eT8dJGkTqT45IavIV
DRVFKi1gr4kZB0jHj6mSdyqW8y/eI/i1HrE9kZoHedqNQJcxIF727ZMnUnmI4OLpYklKhP2UQnmu
A1BaNtVxJ/I8Pm+h93Y3LAihIAYptyf439+9FpKRPY6C650Z5Fccr04fEm0Y1b0W2stoND/h6iwr
4o6CwZqSQ3hee1DVRzZDmtEcBak9cRoGP9nhkdQFB1617uFZq9buY81MYZSDqssnoJSnE2ON7s2M
YfPFtqMzTQsPDPutfcbWyjQ8cD8cJSWU50lMwUpsCzHRFkJVql0jnJdhNlWbIJfB0/RF5c7M2nVs
SywPX1LL1Mq42FrMHGzKayoefCSe7Ha1Si+1PfaScTdLClbl3PzYQCj0cL5pnIOZxkUQqZMwXzIA
wTMklmJS8w3vxB3mrjAh9mPezysWWrAlRXICKGcNx2OXhvJKCY7LQ1w8i5RF806c99Uge43gx0RX
3s8g91qS7dLNXvyEPK7FMbN18OquY/ifBx4lItWubo+TgapFHwKCCtqxm7H+Cyx23vsz55Y9G0o7
upvV6uSCBEWROQKhY4bhIvRnYvahzExu7e+ed6tVyekoUXiQaE3iT+1dxLhIW8gks1glVYbMTzjM
p+lH3+BKyd3dvkJSFF083m7x74eunlkbyW/fbKcUnkuAGACgUSnmR+jQBhlKoOUofq9hmX2P5acc
Fd3juWlwT9V/yo/Lchb2BmOQ8T/tVcN4nsBgbFHAnFeMQsrtY90goCeQ4KANwHoKM0PG7mWTw0UJ
907rctIcLNl2Q3A+FgKf3WZFyRFD1mYVAddOrkARu5NfdmsqJIqesJ+w6toqUh3wdqL6rQxoc1FS
XBV/6S3+17CUzVjJvPhi7FAiuvhrjrfclj6evf8QGfkexmXfp4iNDzBcs8xo3DOf3JPZ1NpVJGBt
E3Y3VKT/h8c0qwIFi+7ArgjTN54XbkfC4JvJZW415JVmisZtvX3TNGx0VsJV0DOB7qwVaob/ii4L
coBqcbyc61YTpR0Lr+J+TeznfdBWWkPJgw5mrMyRYWWHrWEy6FpMPzZ9U8UVf5Fe9bJrPEhjosL2
0Ypk3c6ldPX+izDIa99ME/uy4tQG89Q0y+P0EHz1iwioK8utQ+2AthtNv814lDbecWLE+kHiUwqe
Kx3Ly1PhDcMe41hHqhducxcEfbycLGh+VpH/SDrHH+X0a1Bn5IQxB+GN7rkgZW12Jh3pu5xEq2FZ
B8231VGbHGLJqmUOwRZFE3TiC0v38sDY3M87LwsSnJ46we6Z5Ht+jP8b3NyALE8licLFr1ygGiK8
WSZULsNolUVv7XwnOst/HFURJT05O+rvApjTN1v36C1xBT4D/PaLA8MdRdr+//ATb2n6zF70NLcN
le1bU8zaYfcusHUDuolK1eFzAqFOycX3ICi4F/HsFYXTgL9YPAGVTHAxcIWf/Dl8dacWv59Bh5Db
i+1iNntVMirXd3aI86QkXVFBqSfyXHe4czIQ3LDbniIFdmCtq3U2yqf+fO22Vl3IYZppD+XBYkq/
o23z7p8ZmIsIJ3lwysBbCub95sXy6IhzzgiTz2ZlvJ7i+dkYkpvaocw1m3RmErFgasSw81Hv1Nj8
lx3fOSQmHLliqHuDnKZTVGVZym54MauYCMIhjhgQ/JM9pkhf8yj1lLRuVVA55gGiCVp2JKnu+UMs
2wYJkJDmmb0KNct/ZSJyqjYL/rV2oxESokrd1pW0B7r8dCLmLQCxTGBluFjpxCHIAhjdj1vrLJZT
o6yaY56ufR4hkrXms5tLAR8O8uJdrpho1uh0lc2pFRd8vzUwBAo0CZqed/1/7CRE69z8t0xa7rt7
Le5fHcTTKKDKIPNpl/E79nVgqYEzhI2UopNwkFH9rjZSU6iJ9QOmnNPqiGxK3MchvqbKq6mMj1i6
RQI3xvHv/86OYc7QQBPrvE1pJasQ/mtkihlar3XLd7241PaofgweVWHg1KUNWU8z7mGr9+++9bif
Fs9zJdLCf8y1dPlQhSW65CPxacjM3BljbrwE4l9r6uNF8sKrNBGRUTwBDI0f/6+ipO1kYxGQMVuv
VDgfSRisaP0Tdie49WfrHDI1PNXguJlV3v5PMN9i5kAU3/8+tTCbz7gV2K05uGL38n/gbmMOQTzu
OG+ZrPlVD5TWaXxQKjiQVHt2IXepz6k+ubH3kUiUHCocDFhX0xRUip6NE0IK6b7h8bmtM+hzs9zG
P4SeNoCoxLvUakHZw296NgOyjAhyHgZ9mJSkOBf6UooM5+E+Oh1infFZTO1/4PbkGu2QMYGYlSru
1aQ9QOLlJAYJ1FhrG0fLGUL45uJIotwc81c/lTEoRfujrc36g5iqujjdPP/y2H5VCT4wGNTtxAvO
WPK9szk/inRgUPqmUnNzjZ9Q6w/IxbaydVmYz3NM4cI57G20dU3adZU0Hcu6u+u9Navn7A9I96Y9
jST8dmK/SzpbdYkBxtpwICNLtDl3e+O4eRP231dLOKVLk3fOu9hHJtJT3/7mVKx6oWwCFOtGPu7u
ZxdysNhuRxxhH/riZ6IgADW/6UlLz2eODmtCr+GjiylCbfisXR5JKycsn1m/lJWLIrMaLhTbr06S
tUNXbimu34it5A1wPyszeLJycfpVHLhG1XRnOzcYGKxkSWwju9GbIic01NHxvNwrZCKLTDjbsMf5
BHiwv+DPJXJ7eJlIghaFRk6Ez8Jw0jhVEKQuywdgQ0G/JkGWrsj9w1AFymMBRzCwMw8RyHnyPT25
8uW05uALROzFVYJYpZve2UXGHEDza7VIT0B36/5bUY7bZX/T4SQ72u1dumaSZ57FMzoX99nzRrpS
bX6R5BjChw5Rtc7s1vbrQcmNf2g7V0VEYbx2fCRpqccTGc6KvnI9UfXv/j/5v1kYCbnC4xjqvk4Q
f3t6w2wOEhAzUcAH3wFB5mhG7M5W1kIn3ZL/t+5K7QwZQj372AMBrZcmU5lBLxOEryo42n/548x2
4QeU+bQlLW/d1UP373DOG/QWdLE0FHEOEbvUaSsSatiamN2pXdRv9UYdxgPMenLorSApOQrPgeXF
WAjOdosvuHO73RXp1enu33/5+dvp7ZABkotqBBAR0CVTrKZUJRliIbHQ2mD4b+f6k/436qxHaQCZ
KV+Hda0IU9NQR4Hq0UO0veoQ+By5hcnDtsttowaQ9By+e4f5U/FOx70BT996nHED79Itm/bjitZr
Cu/ZG/0WlKtIh6bjTcIkxrC8fAipzVwCoIj8QIkrjzc80O/9iSk5hx2DwBNxG69HqxfVss5fdJmN
TNB+y4EPIMULfaL0n08y13u6VIYQH6mYqc47xHLLDBV4m2VcT1CsxpMTiyvLHC5+xJ1M9DlCWvlo
pJcgESfq+fn6d/DyIReX5QtlJJVVdJ5tVQP02FPv1zJg+G9VPlYlMRfiGeq9aHEYkidqN9kjYn6P
2SimIs7v5wDuQwjfJxr4QLNdVHRXaluXKnpuIN3TWX5uZhhhdLG7ravIP9Yqbdwv57QhKt5htPQw
bbINQxI4AsWLFBOQJaVsfuxaGctW2fpDFm2P6GiZIihnx5Gkw025qu/BGAa0huOuaiF8/ult0Pj+
DNHmBVCtNXMhUAaDWaQAvvZIyg42hBepc2JiDRePudQop+aXZC+yUkhhN8Ijf/s8sMTcsoYD/cKr
aVzqgDSIKTF/zIQt9OKIybQEuIf3SOTIKr66EwqgnMBB/8SnY5pVNbCur9aI5zu8j+KbG3ZdvTsx
kGp0+VTyE9LD02tTmbxSjABei+XnHjUbIHO2tx7Cq5qwTLBoLra0+z+1QLSKf0uqJxbdvM/ISgnL
d6Tn1XHkeZtI6SgVZVLyTmq/NISXImrCyJfAd7V7jxshu6DxxybQ2M3rIRkAVMCk7NyZyNy/8Eil
khL/ud3DvaRvJsoT1LtZNQTf87mjXtssqKbqABhNGHScNdQKnx1HOhUp7AuVSLB4hyNwuZzxJlEZ
J4+JI9ueQR3bQ/e5leadoeB4lBPy2S9PVJHKY2yEHbCZEVzUTnznRZA2CVZpRZo6Ei70+JevglH4
euEcuikKcHeVZdyNaseAALt4liwbH0OPbrdRKJpJCUjKLi/K+jN8g9qmcy6tDCi+y2PQ87nmjRdq
Ge4CEDNu+Z7gnTbPYbzDINnpGbj0fHEdckUijmiI5tO9B7CjTxziWhx6/r59/wEmtWw14YL7M3JV
FVFeLePLChpd75p+eMSaKpXxrHD8gA8cSS5jKa9b83F+WSwX2XY5LSPeBUniGF0K8ybCHrGmF1uT
GucZ7mnqcAMguqPwoO8oG6+d56Ppby/pbxBqY5sFA2dXdRUIeKfGCCEOeRwt2dO0MuUvrHuCZpMP
T2U84mHf2gxzI9qenLNYAuKVboXsD6Widp6nw0Wnp/qhBzCHNPS/cCD1iMcO3Qy6MGiFNFzr3qx+
3IUNoez5lxuRTkNoHEFgd9IgjNm/eCeS8yl/Ipd4avFSHfG76Uw69GoMMghTLWeN8BbX3q45lPRf
4udtn8J7gIaC+WzDWV396J5zvpP40RO8bOZKunAHeW8hxrlrk8H2ANbOThFYVyzxXY0pw7om0JC8
wOk4QLXVjqbSI/hLsJALDrYqdhYe/lbGUHrGqRuz57qrbyc0Ep9g1lJGecEIhvPREH00nmKqyS+q
hCtxgRoOEXCr1z9r1bhJVkazs3RmI4jgOCq5Z1WqGARR5a5Sdtn5GT1h6EQ7F9x78iui9g7odTpe
/j1VbhYOCxN6ICerkJF7dH5Fp6b4kirmFJqaH7kVF0RUUnWqDFAHLAepdx51X2zRrQtWl0hVk/PI
Ac5/6enruiGMHmKfG4aDdd8rAoNNMqvp0Glf/qxx3wbif7PHp7GHOuGffy1T/uNyd/a2jF+H9Jqx
KhQtFuIBp2d02Uk8gGbRGK6fyds33oa5yZwdFtGPuefswzheg7UOsW1fWeGng/oBGnPFMA2sHfA2
Y5GYeQtiFeBk4Stx+qlgNEcpH5X2KbW+qGLE3q73bvFHk+1SwjTo2b0c2bSqQVKsJyVhjYEhzjhV
s022ocTJaZcF8ZVp/dnp8/7ZhwFDDr2WmHG1BAwwrQZLDdmaNvCkB3tS3d6nRa89aKjN8uIhe9jp
A0M3Mkdp3ZHTLAFqC9i40WnS9pKISrcGHTNWYNlWzoAtqC6rSkZ/EG4nhgGT51Ws6Ey17Vlj1/DK
krnpc+GORH1mzMMOvFQWnh6IHQ+Pe1oloamRUdy5RjcgkxmN0JQOAylDmwElug3GP4jmKKXgK6Hi
o6kiyttVc0w0xHUeX2IBisU5QIRXcSWzMus4CslL2OqgbRtl2ZG8gb3aEEE7/Uqh0WYsRl0ADnTd
bb1XwnQXySBGuIWvXfiAVFhXGn8ehQHsIs7sQMEE6j1tb0qbWxXvSN1BN0Z2/aO9mw3pPEf4KRRl
dWfirVY/raD2BxHaC7xdf0oGlAe25GcBt5Z0zUIQi7w4LprOP1DbA/l2JLDa6ykDcEIeulDcoZCk
0ctg/xBTcBjnECjNF4F/mDwXKLTwyUAhP6hBpkc86XCP9TD7GUs5j4anvXyd1pd2SI06u69yA0ZX
87HvBA5tJQhd718qisGEuRI6d7NR29JwUKYjbUyXNun4VWBp4yPYnDf451HK8z0h6XS+TK2PBWKI
u7Gc4o++juddqx5bQkPFJWHuubdzSWT/A7ue+1Lns2f2FNHMw+BelCDJR/FC5RdY+HdSn7Ut+t3X
/jfnQKfsGBwUb7L9Cj3VXs3SW+Ub7ZdhI1yrD7MA1K4zr3HrM9VVz9IqcgKSYwK0xt8q1GrsI9Pd
LVU7L0XdrfjRP38g9bXQI05Ia6Dr6GIf3YA4R5HhZtU4JFvhcCUpw4GAF1bp5VYD1tOodhw1raCz
vAv26mFi+J+ks4aSk9iAuAh+9aGAPeSaew1N/FVzX1jUsVNYD8CNpT6avsPS7agbaB4Ev1tlqQJS
ufIioRDC2pPA6dYf6qOSTzEO86wZ36YkhcUd0cNCN1i1CEz8zb20KNaNgz0hOunkDoFAClBvwHrM
DuBWcYAnkm+4fbi8SD84Se6vEWGrZjRxilj8bKmTS3H4eTpvwqqSzOc6yqOHM7as5WhwRMK45txN
X1tXHU4btn/A73aAJO8OxSZf44JniN39aLu/FSA6A7JN8fPDI+I4WgneJwdVLbk0hGZu250MuA4g
CryLQedBHQPuuuQ8CyozKRNxByq8MB97I+gG2uzi9nXBHbKH7WY7tVaUWCoie+Iosn53MaMuIY+P
EslAlfLa+Sc0pLtLrFhf2j7afS9q2bY9mkcXYhob2HsUVQPLezwmckG7SkbT/ZBzVn7bhNfQEtWJ
pIrFpIl96u7jtsWDF1cIe7I+EEJaB3qG0FaUygq5jKwu/SazTfDX10Ma/tHta0PiuiV9bC9s1DM5
Gfc5iW2Hyd7/J4pRDSzgfGXNGGqaJZ5KUJZKY6mBIfT3WhjRQ+vboDQef8HUXIhBLNmkxiPWm6cO
PTTJD8dgCi3nKSmu9uXKH5/v+um4cwkZBGPkWlAIsqt88ji1Amy0EsxQeQhngxkrsC+usgYSWRIu
6qMjJBx4U1qiB+1T9GMoKcDIdAU0R95hmTWi51RAAXA1F8Y5WWB7J57EnkVjhzxeDqFxB5a77hkD
Rw1GgAdlAjGFbySav7U5zCNsD+sbo30tOL7WXGFG6DkDDZmpgnAtKG6pH5lekXYDT2aLGAjf04Rw
1/kPhKUozbhn1FQpjUoBeDADa3ouqbOFnlUHXzAYKgN05YhQo1ri2UZxcMBX1/Xv9JdfkfPILbxc
sjhe52ETMZHYxnpGfDDycLe6y7ZttCiQ47SqPty/NQqzBxLiYYvdYkCY/6IwsNqW6AIYTzdatPse
ACLB0i/EG7zqu49Cj09VfqdopB8RHIKIkk6OreuAWJLlSb7qTMRgvVetbtkHIp/XWWbv0QHdse11
XjVIV8t04z2dy8QikQcTOumfnH9+8WT3hhtko8VxVfLRJeSYWtYgYEEyKAtNcjBqRNygy/kJQWXC
DCo4bccoAnC1gQbluhxOxso5mSXCogHtT/rOkXeSjtxnp5y5Cg/Dmnn33lYLNzv92EsSDGjHal2C
CwbCyYJQEu031GfowRAAhNnTtzOeZtkwt8cKR+XAdy0gUe8wkWqBl3g2AzMMnRItpWPl0sI6dlv3
GfAxv0mY9VMAk7O2t4pKYZuaZ/OJFYDnPFZoEWGG3z5dYyejJiv7ynWZH1xfL1iSWb3CAgzy4vu7
O8fkwJjmpxjTBH+2ArMvvdrUsVAXwoToO62wbnHm3Yi5C32tBltvzmwHRyTJBe49h0NQX63DnUx+
EEIrQU2ZYmXPiqvSTgGJtLxLg/teCEUoA/nrJDXdDI3PRhJmYHXZu07/dIK5M6t6+0W1JX+fgqZu
XL+09Ix2qmvo+zUD4j4V2GprygEIDrhSUvCb4HsAYCex0XPt2LtOAdhsc5kK56iipcKAupZP7v5r
SqLAioTEDZBiBFtNmATl4xl+isA4Ed09BbS394nT9xT56kHrHQ1gQO239GRw63NU8pZ/mKQUF3Li
T6eY1lrOkHRq7qpne+ypQaLiiI7K1MzG1QKm+8BGVCHOZN0XsYf/M0JwG5uaY2HKjuEWELSQLnkx
iycXerVqUishRMqQkba97x95vMSXljBcptUl3b2wgYDniGb3u9heP8qofXTXtauD2wRm2De6Aypk
AoWYAV2v97Fi4JTkz/i7YIrk32bO1buCElczQmfv55Sfx5W1B2Zq/VFL6w4X59glgFX2ADvtbNFy
aFiENPn68nVwy+KIyuAH2nTrO42V5vcQ89MWTwckgSoGCnOlZtO01Sgxju46m/SUfZfxJ6vZv2m9
H2xVK5vLPvbb433hXZTLIxT3Qj6PnbYTNk+z9reSR10qTEbPs9aO7Ehdf/qfo5akynnLeZYTw/mK
QFzCuhzOaT4/9y1vSNuUY60LyMKLTYhjR0J20SjyWNcBsfYZRzn5wPAb11fT9MkjdiuAooV4/ejp
Xs75n4Jay0NHma5DHSasgh/YkBLRUrn9XLwBBZFAxTokGd14IQhjhJVBBQhutR6Kk9qHED6dYHPp
YT76MZ2PMywm1Inq05w5cSwiJS/eckiB58Zj1m4RJ8mBsLztvOBqL7gEb1mMLQ5tR6eu/6XdwNY3
wNQ7jajYjvqWSh3NMSs1zDPy2xgbLpsLhWPmklVeAxpYi9Lw7swLg7Se+tF1CKqoIkLxc4k1A+Wv
ErW19fL/IRdK8xkbkACJSAOh3jnZ9X93ty7/I+AvebgU2Xnwp2CmhxnVoMgm2irvVUxVYaN7NcBv
2dt6i25xKRaRW5+bXeeC39yxlKZD7NvpAnzliuQq8lelD60VNEq1V5jkgnjv51NIafnCIvSxlKJW
6ya6p/xDbNw8Ut01eyMIH8errXKja6LIBtgN0X/9rPni2ER8CmxJFIgGfTWgiqMEv2WYtmwjevEc
TmfArKe9xvF3asBKD1S5tPX7DyTMQNlOlHVmyNRPfhaYqckxlAzJpiuRhGi/0HJvamQ0XfDVLEDC
v7S/G0mtXx1IamLU7v9PdelOVxXStDdLjfBRd9AKpxpkclNwcdpG4xHcHIYLsMmim5dmFFWk7CVW
66xa+LDr/jPjDTQry05GCiLe7A0PTpmfrZqEZCGMvPlZHljQPyc98PBFvJxG54gLH0PLAEosS9dQ
PbP9T6gYMtV0JD5sJxLb17A9+/G+fV+B2CZlqZf7wA3GI5xk72eVW+FmgXWLde+MFwjoiip0Wxee
t3rx8zYjssi1SpeB8KLXnm/Ue/31UgblYCV7TGk0sshgVeQXThJweB3eIyRTcnaV0APL/ltf7Yi4
CfUYsPUdB6tQFNeVoE7BG3TXWtQwSnv0LZRNT57kRZ9ruRTcqPFyiZFEjj7z2+QVMvo+NCO3YqPZ
idvTsxrX4xL6ATkTehO5xzlLMEaisVgJY1qJrrR5cPb/5X5xHtzfcJaYR1dxruwQgxSi1QaSJKdI
braJj3VtzfHPUC335aeULJhGVE4KeBcW5VAE7tlrZaW48A7b+IvSCAAyYI68GquHz5ZVUv8ecvdK
5liuhD01CQIIUHufabVYqNxUXnfY1t4Q/FHNGbEcd6r5ht8xgiHxe5eON6jvDN5wpk7C7mNC6Ere
wd6z8T1I9PuDFqmhS+/IkeCT2xAuk4m394y9IIhZf7tE9rGI2CwbQSawM3lNOB29Vgl4r9BM/aVV
gep4gN3sy7stD0vWWK0oplaxiHa5Lb/n9pP6QmfSHiGMJelfjHlz3noTlsdfRoUlq0H+fNnbkfZ5
EsCfbdu/H5EWpkVSljgHyIuVlrI/1E/VIxkVUDRcQNj/Y/gZ7JtRHDiJHzYhOpeliTnRSnWu8l2Q
CmNvHYukwbGU7EqBGv5b/WEiauj38s94FcFbXYFK3Gv9D/yzAL0gw1zLIZ7iImCDejfxFzi5Q9M1
clOoE66EoNMeB+yPruQiP5n5PyJUO1GEP5wZbONw3wJLy7Tld51nNRlf+rQSU08tDYsvwIjcLsYu
KPhy0AqqQ+augW9qvC7qpn+u1iulRIPKp68VPtYjARNv3lkv3hsYOj3q7eUBS13j6EVFYsYPv+uw
TnsYlaXv7/Z8oxj9K5NHsFi4nT2qiG3f/e38bn4Zx0cL+0dmGVN1oGpd9LBs0VO56MiCBaGPPiFD
YH0UrwmHy4KqfNqebY7gV7OADBuxUJKDfSURAz/lod32jUbC212IwFY56IhGAmKg5GNJROs284T9
hMth8M7/7Yl9VuLdRhZwCQMD/L9be1wcY5CPj5ab3LcUuir5WYyEZG9yygfPGdk+IwWWm/rxl51n
moegwDRhWDrGCeWbVgmYUzDdx6oK9a1WjAnUQ7aSrPp0Mx2yTjzmybZUMdf5og5C2jprzwSbKBPw
K/QVqi4c4IjGRY2muNNFUzMYBUZahzCjQQrI7yqm4pvMKvLvgs+7oWV2NdNsoCw8kJE+wpegnNfT
d71SXbg5GO0wlCKDn2DRTsuJQR6S2QjoIqBgt1FTsu5J28SaHYRYY8KDoegU0IokFDBXWDlnzNru
CshQB8V+JU4o6sfWiGSjgGr92jAPLAbqqa4IPx9ql1AecrC3f3xS8LhzthhduISyFZ/XmajPKlWh
NCm1ITcsNHnm3XTejyiTtnVW9e7luMs0mGyKSpUF2vEN+KEFhcg2jfMHvVFsiV8fO73O4KiohsVg
L8nAmuyrcTSNJ1VZCAKrs79mDJhqpaHYNR3JQKNJ0W7WIk5Om0qI0XeGrNlvgq3Wdvh3hzmD+CzO
kxiQXEgGszU9Sj+VVN4szE9ohI90E/gim9v6ZFrqmyInx7JSTGINgeUUY0Uk45suiasE/dNVFZgY
V35o0h+CP04k5A79C7nYFBSTbU7rET9Thvz07hpetdFklwO8Z/OgyFoc0Y3m1ovs69cItxvbDNvA
C4edzgGnjed8SQM3yfau9UDIt4GQirX8KDVzqh5dNabLXxsg0nxD9W60NUkzjb2Ato95gTrd5arY
7gXIglP1gQ/DfIEEgHq32OQ14ABw0AfZdpmYMJ4oKLGH/rDa0b3Y5W6EUxICJhzn0djNb3WgxqmM
/rA5sg04KApnVBGomtPeOIUGQZ+vZnB81NE6xWwElb9fPkwaVES/E4uGZJJyWey72wWxs5U4cJwF
yU6U05tIiJqgey3RVZ31cfzrFgexTdjWxI4K8bwVTTzY9G10E7AhCMiup308UjRruy8LTHg7YvCJ
noliChYr6vjya51HHfFClHBcwzZhZOVNPCGIWaf5Ur3VnF6qXdy0lRCepZBk36wZ0M6UKECNH66/
8uLjkxoSIaszhv8eD6qB238fu8mgcR80PnU8HAIsxoQssOU/utnKJ6xviVIpseLOPtOM7PRKL3DA
mAi/Lx2mpbIetiSE5JYH/Ja7AnlUidM22hDpA9TF7oCY3CBaFCYKIgj6UOX0qxwqh0ZWxehQux6R
74RRbwzq90HvIevENMOCxMDL4nRZAzsMH9RbJZt1Y4mzMuy3HJCtY+zMlOf/SygslN4WGGddVW74
AhEwMN/9hZ5wN20JhCk5NDyVYkiYFwCxyAiVeklBNo/s9tQJnVQiTEsdhSe9wI7zksu2Mc50rgDf
o4X5PYQ+qWdVrXNz7wFc3Z7G8/ORTB7fHg0CmLpIesyuoyq6HdpcVAO//cZjciXXcTF7yQ5ZKj2o
KCEG1JYYy5YYf7S4OoL7n60JFifpAsgLTSAzbU9NT2aJG9jBX0nlY26x89NvT2bTtiC5pIisnhHs
KVOUX1uI9+dbHjWvBKPrr+u1M2xYDmczD/pgf4aRVo0qb4bH5lBQsYJOtjpSUxfCRLq3Sc13Q5+v
YMZy22LiOZ6ELLJWpF2XP7AiMuzJlFTphMd4nSCW3wDmw5zKdONo0BvJ7yWq95RW32pmtjq4T+lQ
Nq10fssu7emnPgEFxcN1tjSe7bhEEKHvaa6mhv7RLzoi1pz55YJ4g0EqDiBFNctjSzfKI3d2qrwm
08K/45J3RBLC9haV576OUd6rpF4E36Li7V0TtmqS5IWW337ZXAbD5krcUQONd6UtPAiHHbw3BBsw
TJ7xsm7An78F8w0uRfLRtO0PiRYI+vvJuNlXZXM3CBTKZDA4JNfSe/geUwgGkv/6E2rZASllh4JT
vy/QI7ibLb5SMmbqhAd3DcGk64Nvc4MOLezzHjhZMxhOqAGxHQ+AbE+5mkFuskaE3cj0qtfXxNAm
4jGiWBZ5kdUpE50Knnu6di+ZfH9OBHGDMriQflwLsuSnXZuaX+ZwlfHyjcaQpoJeVpzZr8smPXWa
PZNVKt6zmlKRjOBvzsIvNPUZuHWiXzIsq8uoKiYJ5rNWZVVj0URthgkfa0B88/CHm/HOJas+cfhk
PcXSpZdZez6DIGlIyvekw8nHvETgjgfQjhbwn20mXHEHsapL+qJTKelJ2IJ480gNMuCAdRYXiLD7
OHnkgdCwnZNUzcDeNLMM2SJglKWIm+H/Uwp5QxGHmV4akmMNjcLKLVxKCMcPcIFsl2ZUJB8qpqia
EGJhphm2/DRsQpBArIpp9NvHxE5NbjTQVjfJ9kjCeU9BqaytMK67hXdUi3OgHppLQkaRa1LRy/o+
k0M+wHbXbI7IB+nyAUARK6sua6l3FFtcCILpTYmva1AY3JXvbLN10kZr1p6HI9WG5SriktmxozAC
m4MhwcYUrfdV1XFFAHWqpuG5x0JC6Cr7OZfmV4v5K0W08hu2KBZYaMfu5krdUeLneSHLg8Ecwqhg
4NavPntGMnd1/7ukGDGPOc533EO5h6fbThM9ESYzxr3AmMqNEUz+HwpYDNqfxVHoN650sK8ubLil
y8UEiSnAm47r23RaldFnMW0sOyQjBXbUaSv6Ohrz60at4zi0En80wU7c3bD2523odL26W3zeKtxy
Qlw5RAnIkppQVrsCVspCRJsmVxERo3U4k/3+unMwtNAKPwNyrdA6so7PJoXojwJsq+gJmvv3a5/+
8cdAnoNxc4NMUUC5vGnVDWgkD2NC0axGWg0vmft4NaJM+YZYN+jtbaAoYyS/qGe4ACWHXrZQx5HJ
UkJfiK5sV4KFAnV1X3ol3aAFAa+/MutgQa8jGAsXWFYUOtITIsIO4NL2nIKBnd/qyuFu5e2rhb42
K4aaj02LrTat/BNZA1txqHLDCM3U99WJZ4vleKMXC7Iq7goxVFHV2bdFHeMtD+ZSJc5Xclf1w5YO
jo+4oPrIQ346WoNBlbsRFBLTTxfqwMEImQulIQ3vSqFIX2qDcSen0ABQhDqNcigzZLzOfSrb/Azx
X0QmRuBRttzMPxmcz9TwxtFhTqpwrc2v8EDAibtKym8yvT+lna6q0s3raFCLlb3ifCB3HpSROtD/
udEwvVDjc9ix0wCr10UEbD34MxtgIBaGtH0whRtFv+yWd4dnqAn3WBsqtfbI5f4AvCyw2Dlv4VyX
kuCvfu+/5boaeX007YmSjW1k14qRDjPkl9W+97rWhYEOfZBgGMLgBplj3+0YUeyH3cb6Er9/RzsL
p3DapQGKpW85zY7L5AvPB8Z6HpSQLBedIOKQltrFzDdULyRAbtEhPFSirz/UFTeQ/596SJUC6bf5
ZJRRhMSXBgccokN2hvAiQ4wUkkEQIfkPmF+J70iGJsp3XMSzl/MvFP3MIa193QFStYGIfD1A4I91
m5KP5KSpYS4B1MFx1df1b6fQaHHkIfSOkFxyTfWS8a1Pqm0Vavr6jhcKJW0JLY2U53HctM/NCt4V
4TGyRxWlvZ4CH2IQ6FECdGbG5XwXk3mF7bu3WRNZSrhGZwrzWoyAe2m/ETKkERSmopUSFWb1ponb
b5SUXePs/eF1v9oQ5DZ35pifxrDuh4VUwGamXMPNUUaBRoDa5bw9jYMf7GpaU2kjX/qnpJ+xSSHH
gPiKb1JgJUyx5MpUBUqIvkPWKtrDXOFbNlKUfSfSPln/AZbzlzfjrYMIWGZWu+TecGZv9PcufCxS
mtyGRL1xHEpSZv3V7fDCVBBZGTsdxc6OoSZSTb9WEQXki+Bp3jClUATJXLXQEK4Z8NO3+sayt6u8
waieNdUzFkonlNyoEnOzfOKBiWIttySyuzNW+cGpuIQk9VGkOaRBKXdh0lvJrZHOHtDcfdxcn+H0
Pg6myJKEta2KYaUvPYrclmyhfFngcTBpMBc9w48L1bCtEgWJyE7/ruUyVh9eECRzzA7u60QPbsCK
Qkj4yoiqqyhKVKJhyJ7nPTeZlaQaaaccdFkYf7WmD9KyvfkwCsrD4/RoC4Ln4haG4Ao38PA7V1Du
0wDeMvGBSbtecKe2fWBx9IyS5gZr45p9wVOOnUbDM2m/d2JE1fEDFPeA3sA2NbdUjMi5YIBf5S+B
pL8AjOXrxrYb/q+xImcSZvEKRRtSPtPrcBb5uyAF+z3UAnKxoGAbYOhMVwGjGZxs8BiJf9k7y7zY
Unn7l+cjlESxacrnPR/NswtAzLPi5vFnj49XQg1pJZbW0G6olw/Tkk7z/kE1Mg5ahCPpBYJ4A9RZ
DZ8Rr2hIeDF36YHCduSTwckpfag/PcG/z8GsN3bawmKAFs2j8p5Q8gnbhpIWEqQ3lmyXW0fjS9Tz
WsZrpVmIQNHOXr3zvyYk4s6aes2fDgaTj9fcK8dnNP6GK7x9tjMTg/GBwp5C7josxPURNu4skt9J
IHADGUz6B/lIcc+JGwn2Kx26ZVEx6G4NuajXMgNt4ij4dYLJ77SjDa9m6h0cjowS1PzZ7MwPTOqW
NLE/wAMEE76/tNq/EV5DljcK8FEn7j7BikC9vbfxwlckBzS0CyHtTsob6FhCaD8ywwQ29uWuo0yu
8O3rA0hEuVndprIgjFt+r53urqOo2sDylEySbIvo0WnW2QbuP13K5lTdGITk5Gvdpjpydo76wjPf
V+PZoTi2EQoqm0Zb0A05uuUfky/SErXYE9ki/F169rtgTAkwFcxUzr0uPeKXIMWO6sJUQdp8JooU
agGStD2zkxQ4un0BDN77QWOjznArHibpMSWqigT18uJmj2OJdmgiWUnkc/yMmP2Mts2vNHLiZym+
RIiFQd4AFabGWO9spWEV+6tfHEM43D7JcfwHBdZQKVSA7Ltf4lq5cj5svM6tcS7gG7GQ9VcnvYzF
62hBOaowwVOw1gc1kBlelH7lYAhv60bAB3Bn88zSVSsPxsW00aPUBYgnDBh5Tq8T0Ym3+pyjfezp
PhYlMyyN4uF457xuy5+3+2GTbuzAb9LdPVNS7/X244ZEkKpTSzANaMInhxAJ1HGAZSyAeEcU+6gT
4D9L/iVhQ976KbuHj7Gf9tZELN0teMd0O9LEH2TeeSYGjcVfR8mCkbxxms6S1pBfrdCVegQumHiV
0r7vVNvqtzx8+pNOwBIZ/WFAt2JjcUirG3DVzes8eqU57XbwaC/LwqdShLJLsQTPQxnqqZxxag3u
P5pfbSU9Q7OJ4jm9Tassc/m6/Z8mSfNES5CbfpjBzJv4BCFEFifadV9rqeB+rVv+wWd6RXbGG+FU
3tfaUjDKLJ1ftMIn8Ylz7/PiQ6UGOb5qAlQSgO5g/5cS49EhEUQfn8fvsDw4WtX4/B7ARuIDCIqz
HnfhWJqPwYxZftdWSCXkeBWwUMC/MFcFjHmJWKSUFIoGLi9UFiD4Wvf6sbhKrz6YBZ6vr6MwRFeX
psRId0FE7RLttLDBIsSRoc+gTe/ovDXyvoRCKZeXIqjiKMWyOXU4V6RRmTq0tJ0tjIbcqq5y8NLt
ga7TyHRbJrzWM5Eaym/hwIxaEbEPtjitNNSapbJXJ0FEhOqWlY6R0B2Vax/wHbNRmck5XmCHg4kn
lkHYyoverx4aXRDpv3ngfnaJB0W/4kHBpOPoxUXQQtkWFq5/FWXmThKlpACXc7OtmJI+7dnkwLQm
/dfWOCdsVpSWX/rRAOEpMq5HP8YZVOALfb+u3k00VldsrP9XrO8ceHwhRb72GlvIaaR05bm6L3kF
b9KBBVfov4XtmyFyvEYV9oHogDn3Sen5kXmrKdblw94ULWzuW2Ge1AsNo/obAlvqMIM2M1tMO2z9
3vxgV65hwwKHN6Q0Q6f1Nvh0vRDIv99uqxO7uDcMlzKWd6ydM1+ud2613UBfhR13fnLJQZtSUGW7
tYas3Ig0btXDm6ELmvHCGSzw+LP6ZgH+H3gmsVgko+vGk1+DtfcyJBTTzmk7CMXENASaMNDGA0nq
AheSEExjlw4jMyAPwS2xFArLcHQeSO7DPNNtOTswQAOJcF9GY2cwukoYfqe8ZVX0r/1jeoA0S8+G
xusJUqvjbY84FsLvq4wThptN/jKClM8YuJk3PSN/LudouH1JPgCvI7RQ/FFvLExuWAVC60ebpO/Y
vsWunvCGUxWWja44iYw6zisVTz37SnH8vbY+1gD10X2PIyw/0ph8VvEhTM+uVXy0EmYTN4u1my/7
JdKmIh9YU1a1F5khIZ2ZnyAGpHf3pc8hhwcmqRPFRcpIV9hjhlY7dV+UnqAfPn6KQVAnUfyHErPI
XrPFg25PlzWmRMRMaRPnJEROrTto67F3jphwd6dbGjdIqcZURRw6r6rMKddN2zvTGb7YzTl7iKT8
02w0NXSiumO4xLcj1qTBb83636b0BTkj+qqPiO7GtppGLu+yRwL4cX4GnTTMOqpWZGvrkBDNs5+R
lI14CMokkk5sx4FiEJbT2LosfdrZUGZKbCMyMfTJZN5acLmhVtY4urAhr/Icw4BrvLOYo0NtWOPA
u/sZqNn2ovm5WixX3x/RV3/qREVa9f5p55/ykOt7NPAdsuVgs09qCZEb/O6c7z7P80tPLvWeBViU
7kL5q18CrxGJk2VOV6K/xAc6FKF2OAB55g6AHZNnVH/l5A4mnXHuibsP+GZfq1bqJqta3c4cFTiM
KwIHL/nWTLYHk9wxeMclrGXa0rol1SiGUs1dUntdEQqnjfGs0BcsHkcP3Lo5JdgtJhj1e9XmH1dW
OGkNRTQaXt5ePyflkbC/flfXvg8qy998vlEJJlPRtMoOPNuevebWeUh/R2X8iLPQEb6Rcqqf76hd
UNiejynX1wE2Zx4PbbSTR7ufmigMVI4NU4WoARUpGAIvoI4ZJKOJNwpPe69swGChYuyX4eRZJNgn
ZsAy7EW0IJRf/LSOx+mqYx27VqODxXO7qdHIXtFuChWhaGRbVIwbeqQailWwgst04qgqn/KA4QXs
yQrBg9oxNQe23OKLmDBu7D2Q1mCgkaqiBAf1RWeyGbcJL9VyiwG6ZslSCafGQgdtRxJnm5AkJGOR
AcvHu0ndVYyQpecGrtv6E4ndg3+TSsTXDlMfd8w9u1qZGX6efh0N6J/ZZCtpZMd3gE3i1pna4Nhj
2vUNHA8aQ1jzVA73AHKQOTvkcMQNaAMUshQ2WWnqlHuemv+XtHZLuZKP5UkbhWWAaQtxw+lHCI76
u9+H7BjRta6jWhby3FheSEojr98hmYGQr2Ia7MIB/SV41tX0lh7Hp1C+laBOJLekWfVrOnGdB4B8
OvZHs8hoYDnsDlXcLNJShKcca8KNEioNCsfta6VyS7YHlIv4bEZcQyzCV2/koaqwNumTleXExsyn
SJC+FEoM4oCSRSFF9v4Ub76/4xHPFEgzirJTpPbMO4dzjhoVdw2S7+ZOJ0yL3wkTpSqvVnpTF+Gn
Nt3Xse79+ZfqT2efLdsMq4PK4FJde2zIvTwUUNjMYKYi0wbd+QSvaIukffcP74FLSeZySFOY+NYm
5DJu7HphKjY+KWYe+9nunQbo2IlJcvFx9BiwxMnQGuqyT/2tnAoJpLvXSmXms8IQnWRK2eM+GFfP
IXTHtZ0fEeTI48dRzLsbWVnPHT40kUyRL7F6YMML4gUcvQsztt0JBHOBpfMiuWtkKRlg+R+Qoez9
QUOEmsWt5k1sIibSkE2k2Kp9RMF/WaCdom3wt+oBsuEqJaQhHDuBd/dZHAfeWzHKh8XXZQgWDM7N
IbQQWYGvmodTxpIPIEqPqgQAWZIFGYECcZSG1jYl4DKpizxIO+UVZVQKqBdEQC9wOvv9L5ySV0NT
2JwpzTjPK1FWu4SM6UPqd4CGNoUmqyuso/7LCch3ky8Uv3U+my2uG9+sMtNue5ZKOkaX6CH9Rqq6
6HwjaCPunc19zRXW2jJE4YySMxpN69Sln+MRpbmy3HvaEC2OU6+s9XPbCGDrSN539iSkn3imyeez
npBH1ufJ8kVPYoTuSo4rQCGCoB2Sn8cFg7MLHg14yB3wPomH4nd4RsFmo0bFd9azlCbj8tg5qvbF
62dPd3+PFU8RwmbU5+HuGVAFIPyv41VSRs+e3/q/xUPtADDQMoBZt8Oa9ZFhI9HeXs02kucMug+I
w1AIaVlVHehLN+B3OVDmMUD7t/Mk3Wn928J6X3trn2zNrW13lWaYFdUgT0nkuiv20d3+I7syylVY
4nlXdMuW13AH1NUCnZq6gEfOZUCyJYRBboEP2Cd0IxW/JytbOKiIUQ3CoLo0zbxg0L3Q7AfolVX7
G+pmEnCCfklGv0BBGdBXW7h87Xfa4AGd0oVBDJxtgAgd2dxCwJ3HblOtwYYyUt0uxKWI4yHy/NeN
vHlUrdxVsMOIebiBd1CnWivJdOpVALmDr/EpXGo4rKaig4Jn7PbuztJc8fM5lAVzpU4UDf+qnRWO
/OB98BXQPoXj5S9Nzsbg3Z2so3p250QXWcwhMr+J4M4qbvEvLkSs+w85sfoin4OW5NbISOPdI+bV
UuIYt3JFxthueYsOiIXEkqvLoZWwuAM69NZ/3bgMHTX3VyjWc4r6hqRVa6Huakf2KewoaajS2Umb
xmF7X1LDBmEjMwGokDUqbomAkyRQdxugyu6S2CJnO/D8KMztlYVgb8rvslxgbGSfLLSJSxn2072r
zmNM1lWFFnOa4EHpcjE73VTJ/2c//dbogXSvbFXkzfoEFpi5wcTXYAz04qpjgdLbm0uGEoVSlqgh
BrOcTcf9w9ncji+218cRvKO9A29Szilc97b0F3ozFeSp4fv+g+cdT412UeaFRB5tVmpBjDKVvVjI
rtd0nqiXfYG3WIv362cFU7Dwkap2nODaM6awp04dwuGqodI7b+VWP6mtCjt25He4Xxri2AGsShAK
14fPg8O0h0J9VciwC69IdHthBbBbhlq4+dgBXFhsJ+3/E5U9nexpl7fEwHH+dKrhFoCm+WwI1bY6
AAKaC/H3LHpG3Is37EA2elmK5/HWCLY9IVQYNeP1+Dr4npHD48z7u+YA8CHVIFlOD3MT1YWlZKzk
Plk4QDrPZbCUgVt0Ms/7Mq93D3kUsKgBFu4VpoXg1T3fa3YICnhiSgevYhggPnXJm4cOj1KE+rvL
TWD0TiQ7mN7v413hlXAn5ZhgOeMVez+Yis/pkwe4tWtv2fNb/CRxRGKL7abJWEdRB6u4e7wfRYF7
6kmx9u7YfNl6JTlPQ6rp9yudOH5zTa3gq4j+EtmqIQPDpo064i1ZWgHrXMUvaY3Yxuxhjg/ElZN0
Bqyqy8TizwoMWlyKpnqEPImoHI5AA87FAHj3lbFKc9V2KSCGdZBC6NQ5qnkMUfk2SZwOZHdzOaZT
UZoR5gtb5WO70B3FT5aA8jjXdToPNvDfNb0KG5o81WHg+w4At7lR7SQmlsLJ6lsWrQPpSax4Y4ZE
hOhItv5hzU5ffPzdB8UzVn6NtCPXq7UJcOBohLD3l9ThaiT1JWfdgwrDmsHw4ev8BnlKp4KSxlbh
jizI0btu3ktuTIWPHx1/kLv+d5OoH0yjE/XxGa8MJN8vj5/ikexVzFPxLxJYN6k7CyNW3utIZoI1
56WJ8a/HbdKpzwoC0JjQtId2MkoHTjHNvQOd5ZWJgIBHC3iCNMWi12sLcFy4kNZ8YldDEnN5bPvm
qZ4JmDzHToQTYPkxp0lfpg+nYnVZU2Gq0Jh45hVg23JLe/NAMr6ACMRD+G11+tFm7+NuGczMPOle
scud54LWHBAWUtWwmrO3oBr84UiXFm4iz8uAMac+Lk7GK2egHFzCOyYnLEHeR+2DiIvoH6kDGUlP
u+7+oi73qbNF2W9cJgXkLwDYbOA0dhtFnr5WGYNJjnxLM1gk5qu+ItyT6hwPRGXu7cKFP40ui4Lg
ds+K8uMYh47e0tggPwuGU6rBQhVxn+GdGiuOdC7Qzo9Etzg6gty7DwusPAjhO3yv5Ly/byEP9shA
vvHaYwCwcDvWSVqmbmMQZT0tVgjmxDae5fcBOoNc0q/XnUqs+A0gIwVe312xgWGzwOnj6ptlnl6l
ZCuyhhN157sBuBPHPIXuitOsbZZ4iYMNsUbs26CQVl0ndKqaj+yKJobE9SeX2bk4ZyqzJGRadOJh
BaYlJGaSbcJA23zeRGIYPagcJ9qf1Sm9OsORjbAzymiEdE8LGWyVVMK4PU+iNUKDFAm/lvA4HyTL
MMIjGjjZI+726zfigwsg5plSYeoA73RmiVtwY2EzGh5gxnZF3UayDvcay3YZblUZXDMUaO8BqcgA
V+Bk2tR7eO/EVEID6C4cedgPn1YDINxiLPj0Eycs+Eqyij3qM8lcEwyMyIl/j78nqAw/rRsFQJlU
m9cpMqvy21MTfHupGZgxyG4M3Qp9Qbf2wcrm1Hi7qS1s0ZeznMFdBDGLk3cNTbT7TCCSOaHVuNng
ebmY8eNyyY4q4/C1RwNyzgGFiQLiedCtRMy9jxZDLStG2gOHzXA2PwQwT8AL+Ljoc9YHTTjx8+K4
mn52k2gIFWSzK9YT5WRtvrdM8H87jHkx+fdpUCLjBmU1QIKyF2duVJrC3Wke0GWhj93sT/Y/f6uq
gcHpBNVgUPdGmp45q2PkARPuag7vfpct+6tmWy2O7/XvJmVFip9v64B1tlPD26eGfLlvVQIHsW3a
Xn9StikNe8HHh4Zon1nD7Ji//UzdkjVcrMhXL+3Lg4VKNSd8B8Zb3uPqL/97j1uhBIYrVo9M/ZQW
qIsEoCxNTEM2bzhmO0c30chPEhoZjDci47wzqgW5EUQe61QSmtxNd/n/MzLRNkxwgEQd0nMyqicp
IlHQ1ByBg7WAZuzZvMdbdJERz8r/iiBve3w1+8rASxILxO/gBAXPfQUtlQymYQMonNNM3MQU5AtF
GfjeoBrNtwAgUyYvLG49sESH8Mg5E0GlvrtzIW82NjT7kzDVGtKsDr+hu1e1HfKPm2UvrQjQV5SA
6TgrsOf/l2UlY6DHo56eHPyTeYSW0TdwrVCy0uFkb0YGAfwL3QnMSBWOCGGuOglclUMqmdIcoklO
mGVJBTrSYlVA4du2TcEJJVvKmyIItt6jvuv1xDi2ADlgZb8t1HtlL9fgX2q/ZoUptZd3D3I7fCKs
01/DV6o20XEGdo/z+V5aXnQasojw1VBxPIwpxJ5N4odZui+gAhmJ0UNRKsdo9nvQM3zcQY5N8X63
7nnu1gyGUSyzoE8zjpynFldkvK6Lj8fdO5Djq8VGslaf8kYNojGnmCYMCh+3bHmObDdfBikn/Qb2
9HdohpQHSyo0YRwBqgNVJF8jbZOL9jitOMwYfPcMHJQ2l124PUtTdwyktD7lqA8zuwSh237xty3J
lz84fdeIqqa6GE+XpT7CyYKoHxMbQeB3TYY+yyitH3Da16a/IDsyaPy4hRXwnJMxQcFJH8IkLJW7
17u5wNKbmSOtiX627r2MFI7SM4D9k5fEPEjc5XNxYPxlCvSeWjm/SbTvi9XvWWgWU1c00cc8BenK
rZW2kmZlkxYX3eNMsA0WKPcH7vas9gQQXHZCHyrV3IlUG5cDWLgBhrRvTCKHuicLCbB4y/7GE++2
xOZWt20/P0sH7bCwP1v6xCHXSW+sFqN3HB7c3R7zSz1k4dEUrKxoa7jy+Ft3c6jiXTkBd1Sqv1/v
IMdlTheZ0m9sF+lP1Gg0Ds+NAOAtuykt1DMUoMAybVnalHvvZ9QbZuPGlkokzL+xFcOz6ihy/6Vq
GhxHhuoRSmFwY2gsKM2xHKYKRuNtvMBJceuoIlUbihr43cQhp3hMq7Ermu7RR/1355NdeU06Y6ML
H78CcHkYmmjvsiS2ESNA7gjEGpLtdQArxPuFvFtjEjMdAkUIxnU+IucKUprZn3KXIyQXw0hv2mGo
FuY8COtlBAqbxlO0Tpr0gYug0a/DuoAUQwqFOFHmv4tWOEeT9jPAe1iBQ2dCTT/NDxKT0RQjdUzN
Pi1BiZ6iF/EB/Uo9Zx1C8foA3hF0yoxW1qSVJDm+9HCY4nUdN0AmmEm5G9S5Lk0PnFDXYNeUQUCR
get24orvDts/gWMK8tO2mPpctV3O0RpkuA2+gBDrYan79zJ3RFD01iNhlD6NPuRAmUtt5ADt5Ftm
g+TyfVHRW6A1U+c1IT7AfMAVRdidSveNUVbB84drpj8IArGNT4QVk3JIArCx2aLoTzUx+EADXWJc
DkMGdRcexCBWgN6ce9p7f23yZPONxmnj4mxAVQD5PAayEy8lbvH5GYO0MKzfwXy+p2KnqC01ntJF
IpveIZXQE8N5KeJPrHc9LoOdCgFEUCqJpRb9BCAxW0hOaD78kA0dqe9HXnrcOcaQWOcGJyRT764l
u8aYZYt6/Sm2gSJls+XOjw4/EX+VHO2HH8pMjfI5bMwALQwnHAb+q1G2Sqb0lt1jiEBa0UpROEEu
8U7ArmMafa/6d2B/kFHXYc85J6i1cJj1gP1VcJgDc60v78gamjMdlZzjeYIVvh8yjBYF6VllQsbv
8l2E5SKvafgtwmVWQTsdzm5JDXQDG7LiQn7KTdXMR8hM7o8nWHHxtI/b6CQT8peUfBkcftFBxwRA
Ucq41PvbWALRlDk4kv0KV/VPUlWv1o1A4QEJrUXDMRzOeZIc45fqNwDbmw8LZdD82ETcjUYbsU6c
eLj7/CPn9q4lgUXpRQBR12KR2qFyjbdMCssDCJPO3X6XWVPAdPmxZm6b/xsstu4oI9U6DPc2s1+e
d0lKXb6JjqdHlncn99huqzwpuTxFCvPR18K2nbcoI9cnlRfi0PJPs9Wd4ZXmSL6eZzdeDcVNfFs1
4Hg7oSo7tfpR5muYVR2mMVcqJ3Gn93SsfGTT/moJfPi2oXTuuajMfTJOyf3Sd8a/1vFMuGOMr5/t
7Y+7rZIUzyQoA64OeL9k+MqxDNGUv3eBrjblVHUHs/np9DpePtjuAnjvBzW3k3n86rEb0R8/zsv3
Pm+fT7n/OSH/wAVuScL7lHyK2xO7uGYpbSBKePvMYCi7ywVFllqRDBtdoxbBIHk3InkVsdvsKnBW
pOBu1iyRbQkHMApMxuo7bbfDc5ELHSlnSwHG3tOz9snO5uo/VkbzlmayBn5FQjOo3CmxLNMFsW5R
0vjZ7YNR2Jmytrtpib7/Jy45BxsUQ/j9NrMSrYT75aSzhodlDCuZvfNgudj8nPPgqGd21eGmzZL1
6UYkcUg0aBtVmAbTGK+LrfnM44aXIfOQw20VoVa6+L178Y02J3p6Hz9vBY16LTpwVugiijff360/
lC/xpYbpRPqldcMNI/awjshja6mXsjeFTtLUGB1Xy6zfEJSG/iFwZfl3laQRi8Cj7KkjafLmvK6g
+UXHnfJIbBRY8APBar0ORmA8s9GUy9HZXsvGqdOkN/HBp5rPpUNYygvxuDaeKbEqQzFIZCn1oaW4
M1HSikjmMRucoPjk1ttPdUyc6OCcvUubP7GbTgnvpG5JhkUEv0nWlP9Utf39GkQlXHiB6RQXg48j
nN9HV9dF7ttveRiakS/nyq+C9MSBgdA5EiFD9/9zVLpBc6eaGuFBtUN/E6VK/kxyNPgNb68LWAEm
f9vdpPSbbBry/RlxTuaRjmikOEwGGBH/q5f/ATR6d58VxdnrOU5rCenTRwA44WNnLuXHJweV0sX6
7Jj8xIEtv07CLmeabLmtQQAoYYt0lJ+kYYNs1chpdcGwlMlovCLTd3qUjmtISxcAF/DCTdB2OSNA
0lqAFyaMcnxlxjEW1Qao21gu8PqKfMB4uE2sflB3yFEZknR8k6/SozbGQCWMTeznr7zDurZneKGg
KIprINqcxCw1xUUMoOO8JbDSlH7TneTqddWZtVPEZHu10ZBMpQjuGfB8lTjJW8b2t6yo+Di6pFWX
KmaVO3yvuy1dWdbAi+Uhj7XhSOMDdi1yTlV7mR+y6PgkllTVzz1RqFTX2YRdZ5ktUtIMJ7J4WP9O
g4fF5tqAejp2CkHHZOkpgv/cxPk/nimTP7j/Oh/RfpMTRQ23fsZCnLXRYW7MAjTV3jX0NBXAMc3N
dLcncgnH9DpJA9gGupTsPrrJ4TbslpAfkW/OPZGnbVKUW0iJwdqdQkiFb+VxTrGT2srfzUmC4JRk
UqZ+0gTbnV3bzCnLXI0wKobu0B2PnGPvy2JVBD7zwnevObkK4AzmC6R2wkEJ09oRzJpQ2oWxGQz1
Bkl9rXR/SO4G8NyWn5rhP5lQ42R0fEZNPkqvj3TE8PE3VqFeZxvyue27T7JL1qd+snBPbtcUk2sQ
Z8z7f0hdCswv9tYNfgUxOxuVlYxey8k2tKzFnbTThBCSeZkjwJYeTDXdMIT8Ki7nAyh92EvHV9oL
+n0Dkai1FZxvYkRSW8+zc72rR6XIySgElNcUqfIlV2w8aVLVRspE38qoRhjbJ03bor8EODHNnVOW
LpPLm82nz0R1OGH/vSHAzVe4eddLIz3padmQoR52MqRQHSQ7BkuPPW+zTepJ585PNjJI4tKLctVI
UJjYWjtS5QK+0uK13cK3O4fpzZn6ydQvg31M4M7eWiOaL9gsp+eDfgijoIHW+YHsKtGkqMuEdgLU
IbMXyRfL4TZWTV6Mb71Inu0Ijcpwj4adHuFICkU7trYkNszWcOqU7+fVQUuwq0Pu5coh+XoInmAO
N5YJRZa7CbmwAOPxQKJmGptKJXT/vNVhXEB7GlKgfCzMzsDSNnqNmcDR/3Fahc9V9lYvWguHCq8g
mQn2aPmWIp5ArZiAZ1cL/s6Ew4EGxaQS2J8YoAyXgQhixaMBOZ7jvNiVZJ2bXLuHh4Fz1aG+ZHQW
c+uJQc/Tyaej9uwsNJFXu1yhIeTSLzi5agwYz6LmXiL7gjgSpzIb1sxjm83R5YM+u1JV2IgN/sjv
ggcPSJ9EeiDhJDCvNBKIojBC/d5iEPl6CrBsYMBS/jdfI7RGnN6axJnOIFvDsEbk1jh5UljeUrmN
1upQEINzmLYuTO1hVyuVduRf7LcCxEk8BKGXgUs17UNeUpH3ZOrGsZ063f5UftypF2wldsJGMYvd
ZSTvf9lLS+FraCTu8Wz/zIRpwff8NfT08I6uAHpl/qe3P/YYmWIloGoFxnfbNK3aDHSC0QB3cc+3
jjQH2pYrPcy2QPE/5lft3xPNBZKDzsk8kVzsrCeDoUJqBI/W7CZ66IW3mdx70e3uduOUOpMhrpDd
GfsosgmhtLCLDKRw8e7PlVbstEPEV/tLFPkw/POt14YA467A7hog54nFW5sPYLGqk8oZ747kG/Xx
ofaMzQfDOep0tm74fI9kW03xvdYPJlRPpMCuKxAtwO2AkrwMcqMZojI5UJkv5U/eaYRNmRsyB+rm
j4b3y23lTO9jl4vzeSSPbNf+FOBFg5seo4k11OyG5k0zJ8/LQ+LClZNoeJL5aMcCgCC+lul2Vn48
l+qhCzhvPRIIv9xYuzTU2dMtm0lSLHi5CXGkxL8uJmdrLiHfg26T53Yvttw/fgzMmMa5uMHZ8OLN
qhyaLeyR6jku8OUGHKQfMCZLauJlmoQqph30a4Qj+YiFRm9OSr20bSWVAc+MPpVa4FwM3X0mpfb9
wfifgliqaZrYSkeCir8k9s5G3vwbcfz5Ff3SX224tLFBoiB+C9VHBQMWN1xyM96+/O68j54PK6O5
iLu1/DkCMxBr99VrlDrBOIfMdLK5SywTsCEVPeiGJVzSBlhiViisvr7s2hC3UNS3JsoA3vJylIf+
qjNJuH3RZPHCkju9y42TAC1/HgCUtyM2p2Hh7DOy9ENV8dlCf/LCq055NuwPmP4N1t58lEICURdJ
PZDXvsRnWOZ+rftYeOPXNVA5oVmsfN15sUd4OOIp6qNSEZxd1fAzgaXaCcxfH2MUKdyJGHa4Uojw
7W9nArFUS+VNqh4J9fzAtQdXRgz6hBYkIla6c8xNWifIRrAcdUQVlzU+0aAxYaSmsUa4A0rbONE4
Zpt4md0bOdVHZsHzngFlzPBcIQrjJC68nzuAUVEm5vo+ecij8BcK3xWOmrhhA2unH5vHlySBIxWD
yNs6NW3Jz8e8wHk68hms6NWBOM2jv7t6llpYJTW4m88eifnNIa0LSZsj8GLtiXDF5Joo1V5dmXjX
U8Ecwlgt4AQYovecVb7R6rndH6To3+m81JJDUPi+l38hlYFiUhdnO3YOpYp6FYY2DCoRMC3DaXWg
ADkbzR9vHFEmDiVSomDxjkD2InGmZbh0ntmIu2VlRzGf8OImKw3oJA8AhYoQvJp2oB7prSSNx9kB
XOA3pMnbI+Ka2rrAXmbd2S0Rks+4WZK8o3j5/lw+xhSHLoFSmh7JcEooTSHMoMcg81/M5+TKe8PV
xqx/8/XdhuejxwF14y4S6rI98JkG+fsvFH9ZSFbdeMOxTeq5yQ+sV817TsbkRA6xvkOAYKRtHBxa
b4LF97WAk9Ltbe6Bz9QB70XXlGU2OHPzUKeQypjwk0PZPqo0cqWGZzxld1JqXFzICTXwPAIrlw3S
p4ZOGW9qdYxwQNt2T3YdzgRyhvHjUIXSL5U3yvzbbW0r8bfIBiuTcACNCy/Xx/M59uea4YxduqVq
/aNlWj14PZrxIiiaJrlUab7y5WG7ylkMiNtL441ZAZRPFttiSWvG863J/0QlqXLTonyFilnUtXTu
gS+oOQEgMuPCpwo/lcLC06+JTT64DvxzKVjNriTRVAU+P48rZZjrv8p5CuYb4Hb9jh8HrnWlVaDp
3yx2R3agVFN8tHDTP6R24u+zgAEgCKdUZA3V/k/P75oE45hZaVAAgq6nfW2ZkKUav//RScQhyNuk
r9LGGI9t65DRn0WTYUJEj6FhYUcYU20kXyYGxtUKQ3/OETqAYv0r1WVXi725F7EnpsA2t6cOJmKu
pxejubF0YZKPjEbofu9uGiP97brZThz/+MGjunAKXuM8DYzxSNqHfmwyIuuHHiEWtiKVvGuVT1xD
L+SoLYaOLrpxGPUAorplE05GQAzAPPZINb70HOoFtRqMOvGqJBfl+dF3B4r4jqzFyeEHlLRWg5v7
UEdS/Wueb0W0ZW6WuAPLXKsuE1Q7ufeBQGJ9C1byzKEriNHKn4TLREiKH93F921ShCouDHv1sS5r
i3bueNmUXvhnZp20YuSbvlO2+B6rUGo84JjPp6dPRXnEoL68B2UxpXqlOsjvX+q2VARMLwTyxBCD
gQ963g9grDq9hokpaLBBEAhts6Ig6C/bdaA3AJcwkluIzaNPboHRqteSgTnC2WoNgZ8U8gB8+TCT
6jGlEZCiBVZAa2MoM5Smq7atE+pVjmFxa5+1/2vx3P1G6incR4EOb9fCVnURC4ZartMZbh4nyDw7
lVz5y+hkVy0iKS62pYqQ6vUcF9OAEkczCGH6Sn1lrNmamhNnr7z5qTVaFtmRCyVFxYEUZ6uuYRF/
ZnbthTaAT2ebLQwuJMCYq6Drs//m8PIgskTRcdpzSE9dOy7hjHAS2leVVcufphDkPrukcXZPlnRA
MUtY/+zQ6sHdHpzvq2DPUG3xHHpaDfc3MC5saLyezgFIwzJnX9Q+cSeW3TuozZoGTsR5uqjjBNaH
bNAt5RQWth3lQ/6xPZUGJD9NGUDP+PsO88lNl/iU0jRAtTPNfUlwpS1BvkfMHpxuInQQAR/V3eBr
cjyOrdIwU/sRC0ztD9fwGhHXpkh4dE6/fddS998D8F8M7PP0bSHSvFRA8+N+lM2J2zZsy6hjCgXs
EIReOB3zkerypE2xjbBWR2MHRxcRau0wX0j01kyf5gLO3iu5+TTQWsng9J2G34HgAobH3Hts2BGA
6VRD8DZ7EJERE1mDjpHQvpaHoPdDO2XVZQsuKzzQTGhWPyEnHY3nQHzwD8rIYYHgmAEAuiRR+/yH
DGulbpKpJ/U8EJ3+9UT3aX1I3QIUhqnZ9IR/sefTubWiNCb+FiLwaNRO+O7gxzNJ1h9E+d50u+uv
WNCxJdKpX7Tzh9F0SO52WegcYDeyxCZ9yBIWxl7FcHNLX2m4IQ/VlgVhF19fiiBXbmMCLSoXxBsG
zs6F6wxrB+9QYisjBgbVfQnG3n5ANW7BPgAPVhsytsCM8Wwka80m6ppjI83eGG//674GFSKHz3fv
EIzY/PyAvzlvD6lcRWjhQayHwCZjk5BqThBBVfQTVJmTdgg341cFrcN93ftO5RzNws93nvHXLexH
grqNPKCGilhSGCAt4puHnnTP9kBIF9P1e+piW1rDQbFvrmi5cpNzcwwtbZfgYw3pS3HamX5IBVTe
LcjcvMuNr28qY5VpmvaC8dyHHCnYFlQ7F2zgPgB2+MX0udBOhUgxLFsvvYvCsdlM7DDuHrr39vWL
iVsaa6iXwtjFDaRpuCFAosHntw/0Y4Qc7rY0ZYMe5JMclkwfTaZObZEX2MeBwcKW1dd1wGK/azB3
R7//1wzLPHJ2fT+seW7qWJyvoo759mGOjP6Bvebw1akLGGHccuqG/buo40Wpb4AiXZtInyeTOQl/
k8CDo8SnlAk7OeQSlj8EHtace1ikbr6T/sSpHsUpwh+d3noCh/lm7WVeCkdvaTUET24NQoXtGXRc
a4UhqT1Upx2MqCSgme/KeePOb0iWFbZ5JS/W8ew4+W6bWuSOEqa+/Lvbu54co9IU+d90xbKd2uCp
h2oR9lfmTzn2nRujZ+TdRIT1y6MygduW3QHNeBYaQDCwG8j2N/DCwAr8Fu3rL8XgEdH2FxyecKNg
IzYSWvPV/AITbJZGxSYJjghJ6d/0UYaelZYEglkAX6Y8iQJlqxCKIjiaiytVyowx/NePIEDTFsWk
OmFvD5bACyQPWIVAK2MJ81TRnvrbvKtP1fRPhOpcSczccQNJCp6e/Cyf0pQxWarQEaFF6atV7VLX
L8Lc0UyxDaVAc8Iv3/K6XvT02VCS9ktGgMzAUXxsaDV5F8uAQCBvJZ1nrl0WUXEBUiikh6eA6FfA
p8EeknSCvw9cu222TiuG0owFfsErFvIMXKuxb0f+XYG3JxTIQhbcBOGSqgea8+Xb9ac7a6QgOjnE
pHhz77/mz8qcrq7azDAlgbcyoRLHqipfxt3mBhYD2tEB4I9dHVPABWDseYyIax72a61skgb1KNzX
vdzAXC088OCCUJ/90mOOU28zQk1VbRFRWC/fJXiY27etJOZcUm/R2b+0n5wXP4GlFWlcelLh2GY/
YQNJLyyaM3dfIugf2hmCLx1ZNNDXC8A534VgNd7Qxt8IRWTGdaddWaE6iROgo55EEDnNr+i6DwqM
WDJHYNWH9Qg550hNAlQLLjypjRoePlJSTUFShgQp9yogxvtM3KCAqdtLVKwb6SsjlfGZTs3sg3Vf
pHhqFok9Tb8Urq87KC7byXSii0pTy7Vdm9Cp1cIX+cxtX6QM58pY9jJyaU7onpRZGmF6p1QMDWKd
BY4FVrn9V9sDtcld/tT5Ah8U/zSbItxkpRjtJxRirqnhtQNNwDxc4251pS/jsTIpQKV1jVlmat2b
wjMA7L2NhkJrJc9Gxj0/g4NoS7vbIsbULEeVN//KxHTo79jDLtGNu6xWvnbKA4hWTrZuNTF+hmuj
BfLAcx4sPgKbCCCQF8JJl4jP7kOPFtmUc2bLwwcu5EaMlZe2HIA6OCe+ufLwvIBYZsg5+Jg3GgYM
c+47JIfOZx+a7Yx/vPHcKE/CzwIL1TVQ1bdf0zNMN2YRSOKmhK8xNC1x2dlCzXYO41Mqg6HRv7tj
0/Alus9zNHKY7d9irO5PFRYvjKxzEVnV29cMl7GA4HjqwnNzITwbEmdL1BN7p1lOsxcL58F/WNxt
g1t77FIDb00TcfrzZrbKKFVMATneUtksqlSZvsNClyjoVmedWVen35vK2sDOiOjA1QnFPE29xi5S
anG+tPS5LfZsWAa+/PJhTIRUdj5W3fHBtUJxNKLZCtv3HgM4nxLocAdi7U//YZOhftzs0Pqdq8Ce
NF6B88QCqRjXIfU7Q8Cmyvg6vPOR8pNyqNqwArxIwJSpjnk2WAMSq/gMQ+/as5GKGLlJLjQmPha8
nshCkvtQdd2Ed8DLzQfX91k1MuNqB9GxH07WbTskfqB/FnbqdmHgWXw0ioZfpSLKqADKlO+qxzvt
E8bLttQ+6frgA1q6bITljMW5Z+Qp78OiH6saB8bqiOgAbeQ5LiXu9NdPXuesg5myWcBrUvooxDM0
aVras2xL3isBzoy54fkDNAf3i6evEnkFyxFQowKbG31T2Klc+CsO1dL/NErYSA2pmsediQ2fnzY1
YxS1Io1fIsPFGok14GTJaXeBIUyydhJIwJ4FSmOA0/CbRiqWEBtIjj0E3T6cdU4u+cLZwHrNisOf
8Nh51bKyBdlBZCcLyEYdG7oZXZMGAEOTg1BZbybRReTpZ1UEJGi/JCcdzsyNNmiH+x3LHFMkhkqM
vjjgU0QxhSnY7zA0sRr1c2W25YvNj0QsMq4ThnU+tnYSiEChtwwxNUUjij4ZEoNirAXxuFMSILX3
a6NwB00YCsZAfrWrSGlVG7KqinOG1EXRvC7jo9k3B1ZiI8rqVW0x7VrnRK54GSHGBgrkYfZfALXy
yOUzcyeYmj+FC2D3lFKHWSgZsZg2BlgGZh5VOqqxOO+P9nHcYXT0GKHPueQ4Ef8Z3herp01JdJNQ
nGZ6iOjxq87hPQHzbzmQkopAkWmFHpBCW0YPvhtZIjShJoVhIZ8h5mTjVTvpio8LU1c6EsPKgMwm
SRykWdITCZp9Lcv11bA2Z7oE2pSUztKaTa70hiYnndNJScX+gnSuZ++6DcrtjWcWxC57oLQ6Y7p5
xezPbff7I73XhSeO0d3VxhEV6SwuAA+qKAgWjPuLeHcr07F0rahIR7ex4q7NcNIhUC2VAa1wQXou
a1tknsKQWphWVFzjzzEfj6rSlgtWuI1ktfDovN7teKiufb77Im+xv4E87Dl4gWkjxo0KqiaYUK0/
CHhhf5oJBGvWp2bfEUin5mVWeOu1CC0UbNDUXRnOyn3t6KlcEfE84tMW4eVdiZfZvjo/2faY1Fiz
1mf4/M8J4NCluLQUsoKN86TvYNtxWrz5n4HM8bEf8NRe3Ln/+MtdXuCj5CnLNgmLBbeqeUQaTneQ
USmdf9AV6C5GTJYMcTjh737Ly0lsD3Cl0n/VxZkZkFAiRoczyoyKyoFyQwDPkheHwNQILBvr8qDc
x0exTGjAGLYQvScPV+Czq6OQONmCP/FOjdlOfGeGs3ZkMSNSyIl7gP+3rAEIXya/iuTewMrsqlyD
R5Q829JNaNAyfhXvjpGzyw3EjmVxI1Y4p81uvncB3u7Wlp9NV0HVm1ofFtMd330cYEtktizETTVu
iZobb3idgZadbP4eH1vt2z7ey2bR5zQz6dHFpa6uVuQb8BuaqO6LmgQEYJneJRw3IXu0p7cW6rrU
YBz9klsGIAcbZ4tPA3joy0/1XCptpAxrCWxJTRpw+4lC/LAaWmwvLLm3fS9EBwKQ1c2gykMJ4i11
v0P424H9PwdB5jrnUZdEQD4WaElN1h2xVa2Y+teAXrX6ovBCbUz9xktBNbQBag4sQ4uHewNSs6Tx
0hSvmBi04MoQxz5/w3/a6pv4fHT54h0JcHWjR28D64PAiWVeoLZzx/+Qd3Y4D2FFU2vURc+9jWca
TFAtmV2fr26dDcBVgNkIWP75Yphdk/Eak/UhqZhF1y8TQV+AmeogpQzTAhjgFt3WlYGfDTaIOjAk
aVpJ3ZdVZFLQsFadrwBwicFkQvEgzxdgnzhZnpyMOnpMY/Hulv3VfAsULp6YD7yc/U8L+Xxeqkip
3qbNN08/uEX+8UoYkokZOL7eGxz7oNjGVsCP3qp9P0QuO/o5mgtaXN0icCmbi+uZuNJlav46x7pL
7ShvrjwQLGJXpLzXruU/7z8Afaiwx2VukjbwTk0KArKu5ZEprHFib5QxB5PGl2hxtz1SwENG6qVp
hwoXH0SslhQVZyajdj70EP1oLOGN79enNsMpY9nXj6gaWlruTmSei//f1wawZ7Vj+FOBEoGs+pa6
OBSi1NM15bwlKUCbjTe1GP/YGrlkQ1yUeNVmeR8QTFbtDxfz+2SM8+4BeNSgND0u32T0rS/bVY3x
08/N2URn/VTrS9Y1H+SzuyPdq9ZYacbk07m5d8ThpeYFOX/N2V2r/OR2J0D5p6bwID2UWlwN6cTk
riYjpb/2Y8VgX9jJeMgCf/cD4YUMBcMUxUY4Zp8P4x2Zylau2PpkutzQrPxXPmhHzbCXAVqUp/1r
n0f14NUOMgCGkgGC26exD/cHYLzDsUcKT+6doYnvnpF/mVO6DxYmr3kxGl5pLYmfei+M5ubcW2yf
rzKiD6j+vytyhDemrVa8Fo+ufywpRalOXYI4Htm5Zk+Gx/C1x6OBFvagM7PIb4s+BWHUeyV+BAZP
QWmRUv7ZdkPZDtlprjtR5jq0AR4UyrKAaoItH7cd5Kx93sTZZSkZ70QCwgjcaBb4cigp6O2invrT
ziolNb5WNFZ+32o7IIrm+egfXYGthP+sfxb4Ti/tqz0qD86ZsCEqug77VV47ZbUThD+SkmCeTojo
A6GrMP1em+gEPzvjPxJtOvXOT+fIFTJ7PQ7M94VRgyedYWavqpvFQpAVXKpYDmJEBdYe/9TTvK3l
1Acz8w27iSgd8a+BoxowOTt+WGSxJU8INBiL//3KLywD790iiYn3nUCk4KH0DvKxxw1iVQxmzgrs
Q+dvRKmWOKX6LUWHq6cColL3GL7CuvZ4SaILqh4lK+MIcR4VemvX7DuSLSfl+4HiMD+MxnvcrivI
qC9NV/kRZ+zzQVpLkEd2ZEShV0e3EuBPtXW6IsHvvcy93+x6nURWAtJ3lHrSjepnRuccRHlE9jiK
Yqlp3tiLkEJDuGIkXYhm8C82fKbIS3Wz5wMYQIBTXxh7VR2Q8bwd4HlD9XU8WRq3zWTxqO6K9FBr
dT4xt9o33SarZbq2pIfs6jJiojcm6MW3HQ9LRungIXMynbv/+Siqs0/6tCcr1FFVpqjTpTXk/KV0
XKxomFkTGgnXEc6zJY+emsKWUWi436YqKr11UjLfbXAFO0NhjO/Zfod5WWCMmR68CXc2DQdHhN4Y
VDjT58rLd+zBQU6JdBEMnwZ7CvkvLrPuZNLEx4VlvJCTgJFpKJwkhxB4anfRaFlBaKr66sTZHsh/
8BJlLyoTLRUB2c/bTnXIqKTsnrvPNS1/kYZlyPNndFdeiiqgqGkcSO7jbaO4e3U6G1i/8uiZh1QE
a74LVCTs7o9e33QxsqDuOnRA0nENJX6Ea+ZR8taVfLqr6P2lqhZfbf4Zsxy5nzFi0EOiksFOTva7
5cuH36/+91cW0XzLrne/ouwgg2L/jaU+08RY19/ppm5vawpg3KPQZv0HpE36pfVce7aN4POyQy5r
E+IJBg3F+tE4oaBIM4Vr0CfneQjPrbWc63Z11wy+BgS+D2vMXpv9V+D+B62RX0MrMnwbK3N6uuqf
Eab8YshyvjNFbVJ6jyE4vlnvbArJRaucX1uPhu+04biUof/SMPFWCRWLcM5JNWaFjDnBSxrzM1Nd
8CoKme7XoRnCUh8mGfoE+s88bgB/KunzOWX7hHnSFp+v5New5lOso+65HjL5UOlZxl45e6Yo4lWu
AY3U6q8h0M+8SgWy+HoqDfy+UuzX+tEDopApUlpmqmXvWX0zyvJ5tyNRxQ2xu8yBPU7wLzLW52Vd
rdqYrKeXAeUBP9xfEjZYA4tBt0eCqQKeLdzCUmAWnQjSSQG5LNoNcgV+V21BRcqH65hquEHj5LqP
KRirzrkF6A1clv5fXF31la03N0mKk4hz5jCn+XupgSx4WfulvxLJgDinABfwd078/xZPeUEAAwId
ZQ1CrbzTu0dMDDV2++LdNFn+FJIT7A+jwlgApMETNrpJaUFWnSwkjqeg2Fy8lYDiRA01ugsDvhEd
fLthBgvRXaFDHTHw2isqmBmr153RNY5j99M0IbwZ2bFkGzljMhbWSupvlyjCnOisiL3NS9CQ0zxs
95McTD2nZDsn4AAs+ch65HeuLNWHWDvHQc7k8PZQLZj+lzeomru+Q8FfQ0esBlpyBTHXuxSS/qfz
aLsjQE37fsWN7ViZlAueXcVYm12exaHBcbrv9eEPIvFnvxD4NeSfyg1r7O14TpzUBLHcCQfYC3lM
v0gD/fan2rfJjWAx5Rs5VkH2p1Y+3c4baJY2IRYmaXQzwJoRBG1GzN9txynq3xDJfUXNtI44g8gV
d24pb8ceC99h0GAVbVdnR7kHoclYgGm00C8TS8pqqkKTgkt0elVbabJRb/v8T8ZxiPhWYA3LYB22
sILJQwD+tQ0pIvLOlJkCWjIIQ4FWHv4OjmIpc9lfPkim1mjKs52aw1Y13l0+ONz08GaS+46yyEmW
boIQIPdnFdwwMYydizYyKXQ9LhtaEcCKULFIsZDT3iPyEIWczxH1j4PnsIxeMD6Aj+/oYqN15FEM
0UTXl7R+tkkIg10hxifibG2dGt7bvzEjggfvLE/nyhDpl65Yeq1tvzJi6zJdw+5UeeZ0ED0ZpJEe
e0WxwuQtzjxBJcwn6xuaMLRoAz2Ju+NhohwsjGu0yhegWGiv6Cx9eA5QGV0LkC6bSOMBl24ocG8p
rf+A8RI8ZXtENniMtGYymRXnHjlxFqEJfiEmDNDzyGA6E1/cFj6lJ98KS0daEYPZZFxSLaSMTpwW
IEgC2g/JH6SpUuvfn5QINXIcCc9P8DKg1k7Pw9CFWxk2Ppexkkh31N6XJXTsQ3KarnaYnN1FedfS
jApis8QjWfAoZ4O9xh9rdHk1TD8uwGpS+neuurW42u9MqnjZ2NXw1RGzceLbWFbgqQl48rTYv31a
QU3faeV3Cqt6rzg89H4mdwJQvKTfYiGrgFLxAYTmh5kQNaJnwKNtBMsJSPa/uE4xj2F40LZWuFjq
HuqaTLWFX0Vds15vekyPaUcfPlCbqNzI9OvF7LUeOsA6gtZMiZU4pYB8fGAjaO3j3D00k/pHTIEG
+h6gVk75yCmI/1G6lC9789qnXQ2FQ8/anxyceX+37ljcO3eUEwGoV9SpZVCJIfugakppo+qIPTOT
DSkz4qtZroxNC35dcI78mMU89kcibH16Pp8gmKEoyvhlOw14yIIAyIVAdb4F5Ue/0S2SIgv0bFbk
L5BSgOMpMf/dMo+acKT8yijTixfymu+1HN90rs/4EAjVYBIWOoQBnB1weM1bmjuFpshEOU5z4Lxn
SaXBmdOt+06Jg1SMoFcRdMWWIQ4ag84SiTfIrwdZvVQihDKSXQl6j29go0c0woSK8HSUygtWKZMf
54JOrfkFsEkAC5oA/+f91b7C2QzgfWmDrGOtzNRXve3fjmPBHERjF1B1zAlDylGseS8sioDUtdtT
4yRmOI/19cDF3e0XmiSP9mX+XHVEKNxRstNG8vxrEqtPNTDW3vMxD4QfNWD6cvNGT/UbneNtMrwm
OpV/2lVkQUIupzQFoj8lUySOoqc3vJHk3RYOZDrttsJH4ouKtx0rAyBLUu0pno3GOpaK6HGSR/bw
tH1TcRTa8cfttq0y6N7aZ4NX1dVBfIdlOpjNhLG31mCcDoP7pjepSzpVqMN+b0IH0tDv1jxOOdE3
FXm/3VBmkssGbZ2VJMTn4hDgPcY4w+QMDu2Pz/4FNoVnk0NkyWNi1/inNf8CLWEpLwdx4tRAI566
PWM2/DV+Sdmqv+TN2Op4N0V/ZPeQ431t37zwAO0fi9s7CpmMjuHCDJwNTmZxdPiTukOI/UeOU0id
h608oVPNlLMHgga0+j3HpttPMqRkCdw5Fyn9XKLYQdHOICx2NEhuNvk8isBrIUBX9wIlE8QPA7mt
UVC+rpghNzn4dgKi5+VnAp604u5yMp4GyuSmojXf7XdbB+z5LvJPen1r53c/Dcy+OdoD+OaDu8hW
BiheaaJZf0NDTJPg1AdDd/GqMPVtYuYJHkalz/EZ4Bn9L7P+PFFX+dgdRFnu2HzhyqIKk35g+gSx
3pG5C4y5TlNooffYsbVIETrIDhGXaF6MrM8kK+q8nG3c6DYWaY5jqqe005/ax6fJVFJhz21BSWYG
bsUjhart0brHilb/7UE6kRNW0niNByTrcNGU0vJej8mku7U1OFV2itAt8JazDZfc/3llHsimMf6Y
8ShupCN0jLyb3bT8/gNijMjUzvTaz+1bDVjcu+rfSacc7stEL5hw0nXo/qRNHncx3KML/qIEpZ38
ImGOadkWsrDog2aU0jvhmsc8vixU2gFvJuZR2STlTsCTemcmTe7Jzf3awz3pan4ecLh1fDsVr0zv
fElFf0nsOvHPv0/RXIhMhw33YFXzwCx8VmuLUVWT6goCsU6K8BhyNuCmLql1zIgQEr7Yqk42Rhq2
xdDcm7xK3px1IljQPAt64s76LcHOmsiBKgz3kHYqbKXWiPz0twe609PGESI2GECrBO28vIER5OcP
Fv2dRvxE7KFO8RNihnGM20ZR0t8SQb10oJW2LL9UZexuAt1AwHNzyCrocxx6OgWe5+L/A3XvP57C
Y7QffIh/huNX/ED12YWOIYDrGJYkpY+5sM+/PntWO6FXBCd/3/junWaL950L7Y3fnSMIUPYrMTpt
YLTfhyaRGAes6M7lbzjxi1HaHG4MXlMchE3QL1gQ7DdB+V4cHDXXQ2d4YpJps/PgYQ8sMyMNMok+
v/k8M6liXWnBEA1WAWlvK5YulhOKvdtC9x4Sv9haeFcjDwNXoa5wEi/cO2xMOsIAY/ZwG7Ii4n6B
0MaCfGCxeRtOkGqbdfXBedJHrygfpHH8h+FmR/bR/PA9UukNz6ezn+ApNk6OCaeWRMPv2HOzKea5
IJ+NORcWt0jsYY/6bGQodzwa3d9d46bM2W62E37H6qlAfDAQ8RJB9JVY9DOozdQLKEZRaCyfTxsK
E0w8gYtEiQ/vxMNbEsM2R4KmbOUjlewvIeWeX2cy0OgEYbLHYHmXenJWvrykqqIBl9kE2OubFubv
pKose+BvGG93vaEhj2mPioO7clqrGzBKPZuIIifLy4zPnE2LU6//dm0lQAu9n1ce5MQIxxRYdJPx
klArUWZGJK1IWsmrt4wrjHCfLpMGcJNJD0p2pMcxyzG0LBasI4ax1DdWetzQN7pK+HJrCiA7ShXc
moQjiaWSCT+iTVUJDPVQJbrjPAu5MPZwhMt1HXG7ezkEJNyqUpY825Vo21pqihWs6eOR/Zpj7ChI
ph3fLKvpjYw6vwGIA2NS/GgmB8qBl1YERd14FLISp8qEx1bISw+smGtMYVfay2edpnMjV1Nt0ORG
Gz7VdQeCjddSbEHZgrtqnxG4DyhOsciJd30xEIzE8BDJUn4rofHsddgorp2HLymKsCo5a3Ogcrjr
1wjeu0QiJudgVNPdXwTX3n6mJBh5qJ73NyraY7xC7ZJCBbWsi0FJQ3zvbtvkvxz3zOapxDAyjc4J
0jjN5dY0LV1YQVwbcYAb3emzpephQEbBypseAQ2aF5fJuGMhXgANnncw8ebaIh7lz3cejjLKe8h6
lCnyENSXU4T1OsRqwlMBu3r/6qbp9OlLOpLLFTlkZR8UoyTPWn3CWSkugr5sa2QdYUhd6duyKTh0
1RUB51QA0U2hSXYAgLE312CxqeMI9CwGFfOUsNF6+d9n+MGOWqd5dHjx7QgvcqsannPDEuHKhgAs
TFZR+BXn9oGROivTHpRFve8MKHYYtMb41YXDMYN3OHPwE/y8JuHtFF8PLbX84xalcp93FWsumEl0
eK4X3NAnUweVREpSxLOcy6yqzRGa4HxkPh44GH/LprfjWM09FgXRpE1NP3yWzRcNUTz3zDWlUJWU
LeMVFbrmvcnhwcNx7hcVFTQvnA7hGmxrMnovEazovZkOaq1yFpUYfw8rd2uxuOHL81sBKpLvBwZq
4f/QCpSbJLo4mGIOIwz7HbcYuIQmSYYcKcI+wd2F0Gjx6GkcFzl/l7hWziHWAGnvw9wtP1IvLTAj
CaqI+amnWmMOiGPUHK6eoTwS9I9Dq82UFnzoBv+bjrQeLk0FuiaJLEUp9o/Frd5olZo7YPQ//qxn
/wMG4N4wH2zLHSvjnghnALo6b52AjFjrfj6JDylgTvVYgL1YWZGeKVETvMjnoA4z25e9fZmICkut
cejThryIKiLTaLvVpaQR+D3qtyh8uFcb1ei+y52xAzRAI//EXojv/+dVUQamhwd2znW/rPqpteq2
JY7fGQ/krFch9JFeqTfScyj3B9D4GahwRkiHEkHsuiArLRGWd+STjL3AobBsofVcAuZHHaTrHkmM
oIRR1Px0PcuEernVS5NaEsSmmbxhUzKCdZKMiSBftHA9BtJ3NKW+j5Zebe1hhrbAJamwJI5ciC07
Zycz/I5uHbQkhR7pBCUOro0mwjd1l5TzUffib8G1046N4GjEut1FRmCu50+hUkYPiCPdcRFSYAxy
JNfdNt07uDWk5bTUr6nj6x7XcgXb0StDoVqS0f/wnyp7aiEBHnWD3tFLktfjWwcGM3n3M9H8mAFl
SIbKq3sMpjPikMTXT5EuoMsMRb7P/9yNj2GUDAq709/qp1kO2Obrpzx6no7co3RKAHVUb0JISh1f
mFuc/dP+Dkx8ordbZ3D1kvrCxuJ6TUUlly2KuTIRLmh0I6g95c8T4XMKYgalB1cy+LEH5DbbX70S
4tHJYQpe97jN2a3HUqLczWyT4wdXqJkDJr5NQuzQpwdHh8BgX/g8IJKYAUgs1rxeumYnNm7Y4kyK
5Mq4eEPnlzlr+i4Qk22WeQq1f0aJo64yMiEIzDFHdfAShMSd75TKKZMSykYZK2p1zDDplMVp6GeA
SiGWiLZlLHdhSiFL3sV7p00DYKQrOx70pbtoKBpxQlgNJq99pxBxpmPQeGrOgab2cFB7BlLumzXE
GlMSsDIr6XtlqAPsHk8s8bBdwd6N9qa/0XAVXvWUpCwUG1CGirfCKvzV6Gj/qULE26uX4UsyMtsx
MYW72mw1qftnjRfAoxUzXV8LKidnwFLoMEk7WoL6EnYlNah0DtmNZy3rHn0hKco7572g4577TJzC
AyqWMLFhAK7nR6CJ4rmqKKsE0ys5w0wyPmrOEqUBy8kz7daFaG8uskI7OKHWm0bs6bACmnXji63F
Q1iM3f72/CWHB/iU7GzGTsn4tpdhm2Ku9cAavNGnTaDZ4NYLG80R1x8zI40bIyUSmMn8Ov3IbF3O
SPo4rem8Suew5WG3vqVzMOoaZw62P6dr6C40XluDVWnkai+pE6zMQpCkco5Kdatu85HegavarkxM
iQAEOqLWu2k6nP0y4yoHbnuA4TMNWpInyeOHR054c7QM3ceuABLmnItcWfZuuM8cl5/Jg/nnzyK9
lKybjkUVYvGnljMH1USj1qxeLL2jTkR2K2DWCGdYDf84n4PvqVoEBTYkZyKRu6jJhAEjrHz1XIoQ
aEIqN9NN0xRlYTmzaAsb5BolmxXvaqr1zAC0JOTzaV81Ra27V4ZLlalgHQsLiHNy1YXieIioVTRc
fMi94oyGviyF3eCLz7fxM177spyfu+Ty0QVbd3VaPf6Ji/Ene1waPg1ETT+Q08L1kXiKOnNEnp4Z
vvTKrzUBpKxvKTr8dI4NaQAwh3Zgpv3c3nNioXUAaDwOFwKybJUAp4cTzNYRisCjuRhfjakAx5Tp
WGfQF5vaDDll3h0sSh1jhsJA/hLrUqVkTphLLEbRV0btNV5fPRYlMSSFmWEWaF0GUmJlLQjsQMJb
zqPeVtO+mDeP9D2YLItFgFqTOQpS26B8+MeCaZuQp9lYrXScQloxiko6WXoc/1YdfTNIT2fA2e7F
B1OhgIwTc8pGQnNqmerO/7ST4ReGn7495QcvfSkJ60O55J44foOST6cS80oDNgdJprpXe3Poz7Su
hLib2Z/2tPEPGojmhQvN+87hTiGTrRQD+Ea6ghYrcyVnvyMDfdzNCp+RQEYFSeRy0ZMXjxGzV9DC
KvKXqxlaLyL+P/9RQJWzLikNMCJW2giVXm6F97eRBEimYVueCiPirJvUmCYXTPuLjJ+nmrZt/qyQ
1I51kSuSTJssK/OrUzAyVOQ7OXnUXw6EhGmli33cLS7KUcxfODN212OLVZxs+H353jqM6Xg2SCqg
f+zNiT21rl0Md7u23+J4C6i2E0WYT6sWPu75RWlB7cXMTkrl4ieR5L18SfIv+2hLv9HaM9anc+Sr
FWZma/oD+hJ64zi9u9zX6/V5cR1zXgApKEl2DXUJuGYld84sD/EO68gaacn5o4uFzqXw8+ZuW286
/aAPrmWCL9aeGtClJXXR+bU0PgEDA0s2PPvHd74t61/Dsuv5PqRcCtgYDZmJ+UoTT9lerJkT7vXR
gu2TmIl2mGYqIMMd5dIDZotETMkT9KIF3Df9gKWBAm92KCozJGs7wNkQQA2gs9r/s09l5eb08fuG
MypOwJiEovmlNuSiA66LGP+WZoN91r6wEyL6HkYZXC/p4bA3lMkW2ws9txn1mKGXciYrXTrvPDlj
uU/gb8f8L+GoLDzn6cbhwwGo64vraG5zgP2D1w9LHGVf8f0QaxGWywCGpBbE1OopuFCmORJeqFLN
npSNv2QYZf+pxnd7/FhAcogBglsYtaSMp4XSkTVh58YgOvBdAXoLJ5znnWTgedRzOT65DNtD7oSn
6oFRukujdC4tvsD9Wcd/hKoJO97BbzZ3bCpG3iB6PkRysil0HArPm9C+0/wgwBQFhfYKhuQpVJQu
MP2Lnvemq/0D25e0Nxi540td2dXK72UVIXjmWwMgKWOzLERKXMeNGnO3kja+20O0XuioXINrFjkM
8TAEhit7TP76N3Hi6+6laPiVrupMAgGBILqzfAuCxOMt4/jYMX6pO22B4E0/JUTAnondCff3a0mY
vOjtSh6OO8Xj0F0VyfCXe2BhP2lJVmwS2fPgeKWo2xlfeTh6ZIZDKain0GPxv8IrveMzUvV7jybP
bftKtuLT13bcG1734qtYFhOVI/6PoQUcJaxbHoRvB05mnm4tcUEEpEdNHv7tvDPjxXbXTJRwwzlw
mC2+F1t7HEsbxx7tMci9OCYu3Qo6ofG5+kmjCn7sthCRFI4q1zJO/HA5i4kY3Mch2fdhuL7ECuIl
YqPt+ficnd5GWIq4+Q68+LxumrYnCuU2NJv62w7EjtsVLTKw4zhdm5iIfyAvp64Jo/WeytyEaUa3
nfw2GS8MMScG82LshXCF0YzoAmfXiP60k8trVOLmp72SUvZnCm1p2GDB6dZHI/iWpGxX4NKRNrhL
4fj9yS2RELLXQLiLnSfEdBg2KyQEvvo0AF8WVBVEr7E9xEzEFcHDBz7BsojGvRSR+eNFVn8NhlWN
BeSPdseuS5+WYHcETV2XOOSUf+M9+tGY0p3sxxlhKQEUKDN7nMctlvibCleZbNDKeKALzP6kQ5og
WI/AUtGQtZzLUSnvCkCcpv/zE+1PjOkor9KYbKo0d40bpifb/lBQnH2PQUPjkRHrnyUa0jShSTmE
oN1ZLMOX/Ka6GL3LV9iEPMg6ZxtpeTQvEAlj3ruizq8BBcOm8Am/xGdP09Nll3rSZhk97v3wDYfz
APvhT6E1orNVk4HEHi7O9D2Dxe4H5GTnJb+PyP+aod2KLfG+kmLtSFuwhjDOtEpAra5ok0RG9PQ2
59KgVGOBwmO7i8nSCXHoGzz/FeIEifCCdws5ubzoTI95mKYAXYAT8AIxOHpdkjtB3ORgh63cEphQ
gCNT6+cqegF1dhTh1oxZUwcjsrYmlvg3pOQ2fALc4GxH/BhRcO9O4RFzIktHQ0jMmLgkGTP0nAka
ClkEPh71y/boItkZ744TZWOCb+ssJPgEfaLcX4ao0R7ZFLN5MOwuUUL+9u1RAYOLXc6tsG1sOLPF
l8Ui/r5HZVlPKk6dhTh+l2xQVXy9rd98rKz5NNs2OnBCO1SZPEOBdXZDAODpg2gXlXMNFRBNqk2G
Wt5VVejDAGjjc+mn0i9g520pZ7zTm8hE9VfXML3GcqjT3TGFdYX/8UjrXoL6e4eDR4U2abdsQJhB
0coM7o7lCb/ybaRofZ4VBLIoO1jFjsGLdYz6aXwjXIbVd7J4EwMM5VcxpllBJrQTRWTMBcWSU9Yq
jm6U3lMdhjRhCjAmEKCSZfE/i1ViGT1fI5juV6zUfCM5uBbNpuOUcUvq3xHCPI52QCpJZ8npldke
k43howBHJpSLK5AVh3fcAGOri+7XgqMqdyY0cvllAxu4VMmPpnMQaDZL4tVAmj+4TPnMqIsKJg/D
yGHhBr7kELADFpkYQuBq79yhoK/qEPhnEAOgxiBQ6HaDX0lsiQLjSPpjToQUNPppPwnemQZj4arD
Q1vPpEPiwbzPLqnxRxuWRUqPaeoIvLZq9WlyYXm/OcwNkJ1IOPdYNh1uLxQgN3kE48CYmuUe1NTx
ZBI5mB1Mv7th0SFzSYdTop+tD0bdcJ5ChUk59JUqdWQxjEYczfACs4aVG6X33wArkBi4+xuXT8UI
f0OnC/k5Q5WcEIZ23TJ1OzAwf0iYplVSFgPDWFlxCYrtfoTY1RXgSTUu3Rmu1Cd4e12tucWBX1TL
vE0EKR2OHvHBJjc+tGu7rSX3rCcb7wZE1VF4GkWhPpTFlm64FB6jIOcjAQ3yVp17nnUyTMrqhFPa
Cx4YCBokJprLejaAFkN2l5AyHnuJ7eBWtgw3s/e+kbBfEiSDgffLN61njK1ZINjSXjfoDmfSXLPj
PEiAO4gdY0v3jAGMAEBDPBJ8cZDOua7xOH3eBTrjZ7d2yX+nh9zQSvo8Ghz+GzEtfW9wzT/gHqsn
e/w/NQK+zWHqHwZAXvPzWoaddJD2k6m9J8W2qzfoRwPvInngzJmIC7ZG25iMsE8D0i30+EVWxb4v
k+GBS69KnS5pHn2eHxYGPj3lwj0MZXrDrgwg94wQjZ+lQ2aRJU3Nd8EV6JBh6yvaM+2/6wWyDK2A
yeWOJVWPhznGmG3J42TZirpEo5x8wGXWAnV/+7RLcPkBOjiro7qlTgJ7asky9rQNaefxHE5SWJt7
W2cKp9hUYQbt4FLlgc5mAmocSpkrYjQUt9ZMdlxRZsNNTd28yM9Ao/bb/wPAgNagMpU+9p1dP3e6
IvLcBC1PdOSpZMKUci2vzcUkq04l/s8Qa4dc+hak7493Hj39Q42f0GTgGQrbTgiH53u4yenvRW6L
qWP/z0T/6D1OdyKxy1cdO8WB8Lhss68V06rQhh8JbgHtSa2WXFc7pA2aDmTB4QWSyWzXpBzjIfjb
f5v2FY8r8D/PHRTyKGJwS87jqrBRua53ZI8SM9FFiLpBAVxSqJ1TOaKw/DPoXoupG3v64O/cgW4+
tsfCqxF5MwM59rKtGWyQVBQWIdD6avY5TpBXECaP2i7kaM/R2dmoXKRwmsxyOMUSAeGMBSg+gP/Q
UTQiJTWEUNh65DQS2b+SVxlUZLBnAJ52CjaXoG7WImwy6mGIoT2xKa2n25eopkvklItnSvU8y4kX
RIPTx0+2hP+k6JlliK8jG3QddYU9w8OfJ7v7D+YlA0NFtr/Mm5pI48L5C0PJwhywOSh4Tf1lL8UO
AQIsdQz3oBGi4KuntmDUlLJ2RpnCEuYNPQAbKiz0XZ9me3iA6BeDu5ndzmH/8LF3a47+9LTULKzo
ugrDX28wp3awGKLde8wPSsPlTD7FFvjmK7Hpn3dZNgGavgtgC6NNgM1IvlqcADF2AfYIQYdL6g+w
FGUbKX3MKo6S1f3dsJap8alsGXvTwN7y6pfOM1BoRgzRASWVjcERnUMalu3IBs6SPWTI0QbBbaQC
WscRYs3StjV5YSksyVZe+B/MUq//NADM9+widnKCQTVI9+79e7uIk5K1+HsGVDqgz8xW60TE5Xa9
6OYtbjWNXADH+Mh7ToE731mWa2qN3cZI2gsO1k8LYG9BnAx90aHYGHsHRK4sRT83TmOOLTVAo2Re
Jq0A60s2dcwWXHiWRQOy6zfkqumDYxKMGqxn6yVJk3KV92v2xkse/0NoNOVfjayJqJi0SpymIrGS
EGBipadosq5IO5gGqs3CdMaXCK/e3lMez3fto7tmEJ905JPPArYIAmoZE224c8ymF9t7SCAXyBrS
TO3aHSR2QaakJ1Kek+aWk3QtyEC/xmNj/WLy45GP5/FT3xkNzjaVdpl5XMSV6AHEaxS8ZF/SUlYN
QZ9lMAFVVVatETqH26s0aDjWS+BnBWA5uNITkXpicKfZd4f/bCYOmmh3AZPLdfB/227BSWahfNA1
WZ6pTbpLdgqhklBlu4lvXenz8ecEdJ3vDLRgTSmodb26SOwGTk6VoxsKnQ0zAAicCwOw9GvOt49V
dC+31F3Y6ZqciAaGwjvO4aL4lagPHvcSD3rntGTkpNFz3bg35Ss7A1+1i52L/gbsU8DvpgAKGq5k
/nwzZV8C83nNsvUEYPN0P0uTGyos0QNDC7dQuP7lVEe11Pchx5eKgU8nDwcMOi/MCw2nhqx+hUDE
w7J9vIkX4YIDLNLpzlv2rPorJzGnBGUAruz1PsQH9E/+rkeAb1joIYgRctDEiDlxgJF5mWIu6o+B
Vf20w9JCi/XnVaK5zt7X1bCCDkDNHLQ+xbykCP9cuGvNNWeCyZiCU/l6jaUNEu/S8HI/ogpBnycu
TUTvrht9br5LDyPzEVR/izpTq34tseKGm9eAJ1EvCQElo0mqGdtVzf2qW+ZlrM6LE5dzz5D7SbJq
UZeuJSxm0d3X0GFueMDzkEVsQ5uxP6ptu1BYEsY1DSVhWm3uromI2K06b6ZLxTQqRbB+WxWgb0E7
E9TmB6VWQMIMuBLD7Yd+EaOmSmpmzEjSgh5uDe2CJvgDMXSsTSIx45F5iNIOedI5KmSDJlwVHiKa
QSMxzCrzk1pLsKaQhWIvUlY9br3aaUg2aa+SRTzIkWi0lMBjOZEkElIH5FEyUVaoR3aQkNeOPXU/
m6J0WXESaGfzAmdwJKyv58gmjV2jbnoN3bQuZwI9wQB7JAXoG+Ka+7l6hZXFzyMiD971rL2kmcmO
4ZMf1Ihasjsc5WgePru5mxnarV3quKp1Ki7AZhteNBzKnm9Y5yzNkDsXquoiDXMdKLTvwpGr+EQm
qzNrPd/y3pMSqBCyN3Ne16A7H3rqX7+4/6Uo7GSxp5afLwze+MyS97s0e8CPKIL5531h8/mVKJm4
Fc4SA4jB5THGU7xt/y/WaObio6ZIY+y2IAj1QxSDyS8Bi39aQUx+M9N5ggOtmHWuI6265a7P8gpa
qjW5SaYjryUf97d4ad+HYWaPe/LUJeP2KifqcQFyu2/FKwzZ1Eh3tFkVbDZ6TRrAnmdDp0TE0eGX
1KwgGNfs9wHSQTW41/Yt4AD7mi6fDBGHvoS6MRkvJQAT25wzDQZuhkDuhsQ+X+nnIdUoHpvUx2Wz
q5haGxihHCMQ08WkEg0a4N2seIzeLoeRpQ3B+ceeI8md0M6SznPNWrutL2GrP0XWgB6lAOiOxR9h
Ys06OKFNDPlTdvzMpGOGLbctg1F4pKy0YpXmF1padOnZl52c6N1sHzHgfeR5dTzXdm4QiboGt/H6
dnykI9Y68u4sOREBRBKoKLW0OdedcetAZn5PZkr/Akch4q/VVAiVdb5SsI6WJXE9DFGSTDfwJ3OG
kqDJu6NZwLebzUhrObH3guiaM0GI0wPr7J6Q11ds6O0HQTQ2pCUVjNnBxMv1Sf2Cfz+CW6t+nDoV
zFsg5nC3ZpaWso9PaBTklS2+uJ9lDOWWO/aazaAT8Qg20Cmz11ORGejHYVN6f+FamMQJ7i+Ylmqr
4OJ+ku8jShO5H7nKaf0O9vSfG4AoPB0qJR/mWM8yJvznj3EwRRVKA9XqtoOS9eVK792BCYkIl7Pl
EvecqXyI2G1WVa0aRHFVEcEYfF9lHR5nSPxAhpjM46NdWy7R3XptO8hSJxJHJl4TFHglK1pKOi5N
B/7Qj51kOTY2w/MF0VcqW3BBzeRFLXH65oQxv0y2cv3S5DFfVf+gyRFsZQVfWPQlMiWbFp3r6VA4
Ntn9mQwe6cNVMPfQqEVT+EzyHTbwt4aRz2o33Oy0Npp31Z1Tn0LdVU2+iZpLC2pW0H3diTbfVOVI
Jig7I1qJs8DiaGEAmkD/2n3C9RdMc6MYkDnAdoeggckaqNsHs7VLrhOc8PHJsyB2gP1c6kr0xmYl
49SQc1K+amiTHyxU6MohCCicWqfell3ORdedSzHUeY0FlqTC45SQae7qwtrZoddksvGVDPsZankj
/LeXJS+hcpkbu9MGqHfdkyirPAAySHfr4l3OMzloogqM6DUI0z9FIkYc5BxMXtF9f3qlaJZSPAiY
ryjxARRBVOVN4NnyoITX4xyYSMGzE1pf/xitSIqd9gStat8XOlSXr8sP5TTHvFTLWfI3qQaNy9OV
3KQ/48WkL5HwJiVsOmtOSvNsrcddHLcXUUrtRcGR9WX2mi27KHNzmqmWbkzPyUquiQYbjRbxcQ4i
qnWWCApibw91oF0Mo0qr8Nk3UELuq4IP5ILQWo781FeI8OYjkQfnVQtN976D9RJHck48qiIzyKMl
4R+6URMOjaiRGzg94FHqgWIBIyGehDbrXVlO47enzaTaYZcb+Ll3jCBIA4kf+YEMzlE3B5o8VFTl
nvHLZ9BpHgAfn2gs1AWL/6BXY4dJ1srtBwqTtwRyk+lGrHTj9j/laysD0qMCm/mwdFR0QKF0SvHC
MGi0fNYVg03B7Sn2lQFeS6Y/Gc/7jdqNZ1DXRstsyG2fEVpkzr4cgUr0vfP3tWU5Q01PkZqxEV54
AhHRudhVZaEjgCeHvIuprtlI5t7IPU43Mtfxmudt58TI+/aqyrogztAIq7Yz7DU0fd2JbfH22+0I
9OmGyVIPDz7VulK5WO/eoLskBCduaWDXJ49w/WsgG+wkC2WIXvhKkdejuC9nnejBYG3qAaztWaop
fmk8JYUgG6GfuFuoK4KdCe4WIAAhEW5oZ3HwmwYgsTsVLB+krwpmZ3Ma1aLb0Gs/VelKY7ggckpp
Zmct+Q4xTDIZSKVXqFs0VYFHFnKoCv9Y6B8CcQJAUQLTDG/w2mjLrQlbhXZjbZzovrjejkZSxKFG
Nqpy3WpCjHsKNBmcqF9gYcHeoc14tkw7I4Vy19CS7nLuwu4RsTqm56KY+SrTThzy7YjbCnVraCG6
Wdwq7P3YKgndIVzkQOD+UdMTL97ez6u2QxOlNFAuMJiVpR0ALQ2e3PTjESi31ZyLieEUkkKI5Dfm
Z6LKDdITldu9Gz0byH+8+arDuEWS1vRimGX8KlkVrjh2QpZ1xB3iRHH9ZxD/91qapnd6W7EgWb/8
FeZA3sHFfpbr9125QvyEKlhe2n5wynJCSrlhsiXGTUwXLFcEGDZj7UvDlXqID1VRNHTeHVP9EYit
lgSvRTByi8BuY0WO815mv+GtgDHJiwA49IvrLCwEAIP7HYj2oSR8HN0vsgKxp3cYqer41Jx3GR01
D3XTek7KjPaEaV7BlP/uvvuisKAzUphFd4eeyudQ070F17Ff2pIDrr5kYWU5VBTNBtPOvKGTg851
RdEpww4AOPsqyll5EOi2H9rnjpkgIHRC5MT6EaSVR2isINJzBf9If3cgIv2T5mn1X5W+HHxJYGfL
bdNL0QmlYUbFwlaw/w3c5MxPF7+pF1R5AXG+yQvSga9H8Ivmr+8RlwiBJ2Jtk1wEzoBcPko9IWE6
A3OCj/it6eQPzERSfSpugLO2/5AsexmeswtU4lu53D1sxrN38mOf1pOKP0H65ZHrNqATfVKVKJB/
U/iT89ey5heLA4im5zoWuP3BMwiGDhH1pxbfOlOzpQsQe7iHQo9uBSUbDcrbUz460X+56Cql2Umt
tO6Fm2hyseB0BPBin7QR1QxOxR1UYOSBi0wSGXHeS8ar1EtSl8xXCtzpj2QUTJvTIBB0k8bSwdGG
C1Xx/boOvFL3Y6RLUvgeUNk0SQSsxAFo4mLFlCaaMKuxM0TvWlcQnu/zNZghy4RehECZoE5Ktxd2
vMoJfmfDZlWiRlHrb+HYZis2q137ZfnELYejTJUojY8znZXdKrSN9u56gpRJxU/84GsL3te8+1AC
7txgxCdKEYqAGJadM08AYoHnqHsPnI5LQe0ZmaAw47KH84tvVh99wu2M9gl4rD2Agw79Ba3mfXB5
zFHCTO/jy/X5KpZAPYScPPu3LSkvStfwyjOu65+czlJGZ8AE5pt+qEKPhMYlozvOoDha5KoidiKk
X5yf08vMiw9haEB6XzJcd55Tr8aRjuCsdOa2SbuEqImntkhcC+Y6ECNic9prkTiO+SE5EE4kXXJh
LPZ8Nzed2AXzZphbcT6rFei8tJiNWSJYMnSkMb2syutr22LCtUmPQyP/cYdEmrL4HMSMLPZhHODp
1WgfJy4tG0UPXw4tLVLZHDDCnL20JK6tUc5CMXxU7rqBpOiO1LHWDUpdBt3DBVvzwOuxvEFJRGjC
pZtFSmx1yWvVTK0AQmxha4+itEovoBdDXwQODzYQd5FZpwQ+ovluyZF25mDgWcJunjzLF/dFep6z
yJGoP1jPA8xgqgC4bj0N+Pw7ht77yys53ZZhY1K2ZRq0QS0egazl9QTUKbmElRNprSqnAYI/nmj0
Pl9+gG50HVAJjDoZ/e+ekbrxzFBSBtocPskKaXifqcPW3hZMcOtTrevKEESumSJvdxB8mHajCgeI
35v90Vr9MGVjBTtgjlNw0WsWfUEZ1u8kBQkTSYgPT0iPJGABrB6ptGF2RtcBdPOicO4ertrpejHk
U6WKZvZOqifXF9w3HG9eEmq2ah155H1RwenuutIwA6Q69SaVfR0LVs4OEsWbZyDCWm338m6zOUzx
L2VuyNYM9li8pzDsRDzxAfv4cqdwtO1zBWAtKycu8qK/235+/tR/YOAmOggOg7VsRlu62JDZfY9L
L+GSXIiO0LhujZ5tj7ufI+I977Qb7xhoZBGsILJDe4twVRzHsA8T2aCTcZ2UAwIrlSCrqeRYPrzt
v4KpJP0qcXrL4kpuzXRhMkxk2KLGbibktDZ1OjJqRsRZcJ3K5+gXxc4WoilPb2g+z+H5XKHtGrWV
sO2US88aEyAKcu4LMkgvGaYZn7dumTkO6o+4FpNYaMA87Ou745UY4c8NnMfcJRB99J9J2n8TZkB4
6OWhjY2IvP25xi/zllHK2nhs9Y4xidk+fSmBTZGlKa5e5dPlFO7lw45JvVqqOmobynCfV6zPe2fD
Haz/Qjn145cY+TSrdX/GPjXdyzI4Ze//DM4CWE03TaU6yj7NFrpjLiqChhz/u3tCKgPFNYx4wqSY
+K0jXfCUoe1BhFFw44FgBn4rtCMFBnYxn1IP4ZtMeqWSErdiZZyOx+XLxsZbi/UQnqog1BMcDxuA
7FOI7LdMs53o9HLgMi1xe4PwOR+IgqpySmMKwpPUvWAidBw8FhYTksXq8iW3crYIYTBUI17aiUJv
sCcO4Dqc9jLF23VvXlGiySxTDXbF74N4SgHnq5sOJTA0vt6nQi1mYaJ0Fk7MJOLIJmgTr8hhrRgQ
66Z7IkxEqZMTt44PoDSFLL7F6EanWTgtuML4Zi44m51OErdUe78U/uG0ZrHXDu2XwGhH9mwF//3N
fsh7Slm/Z55e/cmULaa8xtMMEz8UYT3KgmFk+hsa5Fp1FctDrgBceccbB9Wb+hb1uMzc4IDa1UBR
FMB9FJFoRL6bgCUbfCA7n+5ROZ27dLky3txcrEokYtDiO4bTHO4eAFdGV52AqZnAuIE0dz9x/5ye
d+a3eZud2I4kXmpzSAgFzyzwxReLFxqf52tveaxdLi9V2CjiI+3HGdTDNIjPwqC3SE5tsEEqehwf
e8DR4tStvvZV3DeEVZ2yGSA1XvjxGt02fz1MWhlaDTk95rh8RyECwbEbcPZa1OOjLzSAlB+UEeQ2
6+tFhs7XuGRBm81zvMwp22WCEgedBmxHom2amMwUTSltHKYqumUlGlxHJgDw7OX8XmAppxjnrrC0
LVQjrXonmelrYMbEkXk4E6XV+S5Qdcs/jrrNCSUme484hrmTS0QPyfpR0aWffOD50tsdEgteHws/
eeepzHUSdubkVWls+OcEZ+FuSYPxBPdnPtQihI9TA82mPR7T+6uZOe0s7w6lykjwb3QHdtRujppN
kqRSu1aC8DJR2c7FJnQUxxN0SBgouqmWrlW5fdJVt/a0N2PZqGvKJ6hH51D77PpJymuKW1Vs1onC
pt6Pis07BTOYyWhZXD/sME1NHuYqpIxCzRZ3Dj2vLRQDjrxw/+vN5HkwVoJNL1cA8IC48GeFOPXu
HZVqiMEoZ0eALXIOMlQdSRbeFMoOKlk6/V373u3vAgkDD/uZw9fnnCddhS3TCk+g7PaDWeo5fPh+
x1LcTMUCpiRaABHdv03txKVYQOJGAbRabwDqJ15X5/UJCQ9f0uVbd+58B2YXFi7nvUL/8HsjKP6H
erevU/1oTHuIQ3Cwhjnlpl69pl71p1KsK51aN0NBAmW1FSroUT2yUm9MmORu7rr5qRGs6nbjiqyi
jxom3VXxMbz+1XU/2Fh8cYcVzN/54kcv1i4OuJF2tQ66SkMy1VO+btrbSTsO/SOXcz1zcauE2vB/
3oTgjakbjmUbz5jkCZpFvpH9FUUshvAs3Y34NK4/7YTQ0fcAERr2Wl2xBrLGEwY1+LYrnnqo+NND
cbesIR38nrC3VFb52Fd/bOXRMCG93sOeU9DrIUFUlxsFkjsAj/XnwC1SFo7IkRFM2vFnuzDgxjrn
9El3155s3vIVoKhmP2mZw+GCF+ZD4gMFovCPHsKkmzT+TlSDXGuTYW9wuuIhuJ9LQA76IURUNYaI
/ApbXX/Ab63SrdmQpJDbfHKy9j65FAgv/KH17XXNgSXcrEhCffUbJ9d11WCfee7IT6ZUKsZXn94v
bl5rhJkHkvTDNn8Kxb8uBmWxKss7w6YxFh5DtYW3Lat+9QSi6rO5FGl/FNekVllWZFgWH0xhDv8b
4vFJ6pXgi/Fkx3yzPdMpjQ50FvJDPegyOXIFTJ7JgPIkgM3xCLmIEDkiY6jQd83YhwFugHnZ7U9Y
PIsTKsCADRcZRcRBMB0/j9pogj13KWp6qqgOchrEeHVtLVAKgTrogAPgEoFCayyRNhA/OqXIRDZc
DV+Uk8bnASF/HAuxJdDsxPjxMe6yr6R1cvOrQaLQFDcr+vzjPGzxMLb20I6krxivuaQifq5nGsOP
1DEMlXH1vOV5bTkgFh8ASyoqgU+7btFf0Eoc58J70y7vlcs18AcCYXVo3JMW/zVVM0hgVtAb87B1
y7xCXD/PTqm13v3Z0bBesGdg/vi+EHKuddcS65RWvRyN9/McFadovlqhlI0a99PS5/2vw309Ybg9
ABeMBr+7Hc3ooZkTp4iNN9u6GklO7Bca1xa3LsKJCNMftnj7Z5AUmITf+0NKWEpGc0p/Q9bFmi1+
r0SVkEOzs4CzopiJk0pN8oGqt+GJ8W9w6HGCv47jtV10iXPLarBRWlDW9g8qql1jPVRfoXs82me7
og3GCanJxOueQvWXErq36brTrjKh62lclm/XVhvRjKhKbnJLvINHttzsg7AlTicltEdEd4ErM6DW
7tC5SbpkrC3HwWJ1cjmQPJ5DPxCfmfTwdo+qAjPI/SsWD/JwAb3F4kpbgc57Adcd6T+U/dDfQPCK
zCMGkZ9og4n3Tnp6zjiOukb3ycaRpNAWt509lIiJFq462smkddNSwPWZ/KprIc6SRutgeF/+YKW5
UMJA363gux+PMSdCjoRJVZr71olr0CuXro1rdPN9fx9cLHWwSll5EYMcLMAduJYxIz0fYD5XK6Dd
V/3PuX5zL2LHffvsfdn8Rpc7tqNhi5PuJpzZm6YK0/qHmfJWH+nrt51QeUjTjXBKRJ3wXUlD+P3s
49tJt3gHDE3gnhmuWXkCuJ6nv5GOGHMxaO8EYvRZwHTQn0IK4zKEd+nGnBPi3QcQ6Bo8DjtBxBko
ePPdhi5j3XUkGtiO+qKXZ/pE+t7BPRxQwSthpFqc/h4VkBxnlH1PeP/F1or14v79nCoC5yjZWA/A
pslJzsIb22HXes7nyNjDfKwnnffqK1Ak6p+jS3NTLzppqnTLS31kxryXfPmOmqR8atfj4yWDBqvI
sp2IFeVm9TyMmpd8Z5R7R1NRAdkzOKPwzzWQ9h9qQWus6aCvP/AcXE4T8EmMnssgL12C6Q2M5hl3
+NGAGXt0g500OJGT0xW9X3VS5BijyVVZgeCXTxNChY2OL+cgDbnuRSFJr2KJt6nkUIIO+N8XucOr
iVvz2CTVJiAZ4Q1xUngu65HVzBDKYufLUZ/AAimDap5fzdvm9VVd/kn86+DAULgZ8KK+k7jzHTJE
yB1jwBhgpqSO6tpuKCDJ/AyBsg6ng+m1wVnngPHn+to2JdnByrG08XtaAyIZEIH0HAfCBzJ1P8Cs
+b237OGe62nS1Z5A1qoLLiGSVnXTOrqB6FWAw8ZJRda6HuyUejQDfueOiUOjZSG6dBmkn0i1Xir6
o3Ab69aU2GEVoQVehx9wWRyYAfqo2xhfWHqoyyp1D3n+Iwh51yyjbmuwlfU1GGrog+A5kYqL9AsI
CaqcuURqT1mSSKBv3BexUcpJC6s4I9Xsgf7YXaZuiUrmVVZrO3gU7HBJ85Ye6g5LFoJtMXiEqVgk
SaHoYAukmr9L6Ig5bgEZfLRlTJMaWLWWax2RPljEm9962JKhkRpR54hcAFsEBffdD55EDyXKpLeP
6x1NM7nKxWQJkcVy+IS+XOEMUbYvAkZb43odxxzRQLbwxhi8j9BEV7rmL7audWnoHefmWgXNRcmX
mIDnS8DriLhRobRco3J4ZjndQ+E5HUOZz4K8NAVsQ6CLL/Jm0WTJvykkmpDC4jw5QNclPcDm08Vf
bK0jPmRwEtqabdxSx2NViq3iDV55VVSOWRLEze2xr/NrX/XS0B4g8SZ8E5c5WRsV7ZmWyujiP0Yq
dD3mZvuJHYfps92CU/0cK0UGZv1yQR7LtZP7gotyNk7kKLnYsdNN9XsfIbwJbGqtXiPUP3WyeiHw
+HjnoQn/fJMbVm/JETCJ15fiQKTXGq1/f3Vnknqtk1AO8DKB3v8rL73ePoa9PmLufI/+CGb7ALwW
z/3OW/7y/OQgMa0A0pmfpVPozTi9MiYSNDb8/Ab47XtCcebr9QNYeUnv/oszrMJqABJRKXdobUT6
NstFZmSGqQfIkCZTcJUCCFIZHraNmBJD2UjjEyUiv87Kc4W6dnfJynGLVEFrmwdPQAu4PtoY/99b
iL/k8O/NhLfDFwG6JdB9VusnH44J36yBOOk9JlpvALGBrbrwhrojS27cJqEWycRYFGu7Wqv6tGdL
wh0P7AZocKVyi5dXK5nXF0rlDyuxmL7AtdGtMBCiChrg9NncJC2XSlLZNwAIW0q5sYWpWVakspb+
bc6Y/veH+pxoeOjuN+IJA3wI7F8gNGnBN/NhY0clknxTFPyhjdt3CFajPigRf+rVQD1UHSOBFz4M
bXRTO8L/tgukdXZBPHYoRsp7tGeLaaltmjJehxbGOZp8m98SB7840EbmWMeiKa0LYjE3ldCOzu2v
sBvtkRTcS/fasltmieVKycRmyFBlrCspjRn+n3VJl3gG2NQpnonRhFSj+Z2YHx0It3DmM1m+dRUr
BCZlBgAjYbskPAYZZMM/Msz1SKer4ZvqmJ9Sq3YOt87f8uawM5mYsGPSv6i/6j4Zo0AcbN+yYB5c
CzthyAjz6qXhQrn3Xv49LRxu3KxOs9RW3Tn/Si+Ux1WVEgPFjv9qZvv7H9NsBlWtgvMB0fp6basM
XYMucjRM88aWwWFP7YhDC2hIDxiTtE29L1xd31MtTzAZczYWcL7nsZjnCU1Q8adRE6wW1y9AcOot
JtIxDEcvtBJvaW6/cBKlOG3LA8LgwL5+nfvbgYejPWzwlzq2QDiINaoN5f0W3IFl8oVkDYG/JY9w
gq3myDIY7W13vYf4syZ80PefOLW6HhS9pz+Fe4dYzBiwags9F9esUvR7StI0XebMXnQp27gRgjG4
2waiipzjMknefQDKTYWR8NNGdh48ewjinrVMNFycj3DCgYL//toCKOdcjhf5vqsJfOycNhspCaLs
RLK/A9Ww4cx2h6ghruAITkbkGOOSERcgheqLNcHBX98qKEdYq3+OW59Z1yl5vOpg9dv254OfmUr5
GJ8PzbsF11Euq24Hns7Yg71veyFQCvPpenibjI74AmYhl9IizLMdZYIdJnjCzTt8dfCqsvEB7PK5
Sh4dPPUxGb2VLoVJQHRErXKgwLkU9Z7RAPgeOpMW8B++uOkd/kCB98j7wHtx5p1l5K5IIQ1hUBDX
nL/nabyOurqONWXCkCzFpXPZTmyE14cppTSNJ9ljAqFNuhkFcgY7Hi3TNVFbLNwUB/AkvQRB5Ygp
PdpkRG9p4os4ChwVChLsaGDtDCN3jhhivV/T8+qEnf+ACJQTsf+HW9zK5NRnaIqjZoyLZwd8nDMh
5Phom0yEoqj83fyU02e1w8E64G27uoh+B5o9QYNq6lLVlZaLHGCJaqzhrpSi1Fhx+Q/pKSxnHi0R
rmacWpH0yQTure5UKuHc/6geJuMZOac8Sy8XEqUjy4A5T4Cwjk/ZvhhnMD2M3MtmpJy60tGO9wNF
2DRz+Yz94hAUAG/oNCcw5ZD++DPZiTwm2gFmBIHpWBQrNqQDn7qkXmjsRk+rsgQbClIUnBXcXg1a
k55uhxulZrJtP0F8LUGbkHelKqUCi1Xm2rACw1/gmnqNOxD8qcejt/B691Z+Vv6XV9Fcay1PDTpL
qEvvVE5VpAnNY0mOrVR3oFYBsNxQXt6Unw49ZvoBlZoEWv8Yom2frAUoopQN1JBWmvvqC5DgTAaL
2mwm2ofukNukiw7OTiFBC1eDj2i7F7eJVdJMzYufTo7JNMIeVAruUi8K1GdDU7a41tyFFCj0btEz
oG/JOLvGTAHceHO/tbgVepqgZaZHl3iPlbhJRL1GlUX563idOHBm+BEm6rApCSo0dDkbo8pNLW/0
BlJfU4B3Mn+t0dMenOqSMdVjjGU76s0gRZ8R0YsZyC7Dm6xCozulxMeIMS6OzxD/qLdz6D0DTh6m
tgh2neDam5AdgBGxqXQzme8Vu93of++hWIajBXupqGtzxuCYfbdUEs3NFaKt7vqG/84Ewz9FzF2a
5hd4QC6ta9/Ty6l1ll9FR1FhToHMtUUC4f32onfDhsyi8abBzP54TaWmzbY9UO29nVxhkIALaFXV
HKJI0A1/WCUCuoIsAd6UYks2Us+JSivDA9mYeTxH1WaGHks27xHtIHitWWoPVn5JorYafn3Wmx/u
+lliPUwQOokk2NXz5hPtO61hur7K5KqCPkKF6dTXif84aZSGytYqOMpY3p7RzIX3tMtXJDLLpuKT
N+XkSHB9mOsLn6nKR1MaZuJEGg5KicfEW98q9MCNWAwDU8VUMwzLj5siwgRCL8qnuDPOlJYcO47a
A0tvdOcaPZjd9+9QTIE1yT8Vv21Q5PC5MzYeyol9bLDNClGLL9YRZDSmGg1CxQxDoF4jt8p/oDuE
4IXCv+mdDvA1c6jjy3nbmLyu/UQ6yLrH0jiQzS8NYNFmhUGzrxYdaeYy6yacblj+cHGP0S17brQB
0BOLvLZeHV3bkKwgoiF9J1kDgvuGENqphqefsSNRWnd1qVPinmZiFAi3pabFsThvQbrijwqLUrTX
zrewBXroLVTEL+JbpFqs0akYkOdn7CiRMMF+TPWkUTESIgZfTQwyrgFLgWI3OWiCmJW/pqrGArLz
kzHQAN+Go5UmEWOCVxJ8Sw8AKf0I451OoKxlQQysQ/sZuRIgJuU+McKIGjCyLiZGN1K6vmr8MfN5
h14z1a1on0xGC72k34Uymdcs8+B9RPvEFuj4SbVw93WLtXOnedUC9HO+pNhdRlgN0bvltJQEZ3bc
V/Oz0yZ06c8ILw60ZAKVRPmVBOyTMUDobWcSL9nGpuOgN89Rz7L3AYOJS90QpdfQo6jWwnolHGLV
JOyBKLGijqvEuYJd+459tFTt8Ic6Ir/SwpDOFPdg/Q1sVnrHxPK90vdkVkePZ6MpCsslCb26NX0F
JxS6Q+iRusX3LpXwKWLhPe8RcN6Ev5WTVdPZwVQ4aHUQOeRDnivQP2VAqFjVKokMZEALvbN2YJmX
sCPDQnO0zi3boUydCgY2M85H9ej607h9IY2Dv809tZFmfX4uGIyFwSI3OjnOxYuun4djZeQWDLOP
+VrD7xo6k871MlBBGJEvfSZEr07agjEGEaxo77wYjz7IVg6ff2B/3IEqS5Ez37Cr9cPfvUtcT6Su
aiALt6CugcsEtSB4u5IMmlZptIgeenhuaITHtwXGCmRFd3QMigWqnP1wzwJc2sKLkDIYP7A3NA/T
j8bVGC3+Q/q5GnQ9Y32H4RMR3YldXvMoCfiAI01qZKsF8pM4X/CaUABsjSgLXMOG8z+2cg5DSyzt
MOUvpPFkvp5KtHDCUUToYkJx1F6tokeWPX2BF+Ngt4bOy291aEAO2uLLZU1NBJT++L+lEM7slb8J
b0GqhUeBUi0xWPcFhpgRTTFZyP0bg6Ig1fFYRGj8musc3ciSXZKcgJZJ8KWubpGIcCBaDeCCD33D
ZfN40asEz1QeO6wBDQfKPCzbOoZJaQAfshyJ5wgkfzO9husHrU+5A9FvipN+QDaoeGCc4K1xNzGs
lw5g4LyhXYdoI3gfoQCOm0FeqnkWjD8e2hZJbIFz3xY5AxRcpJiSUDoOxCWB2desZ9VnU05g2UXd
KmTGWLDwAc5ghxRaVUUZnYE4cTR2ZNVzuFJ61MjGES2jPIbP4f4pnQN5TcapQpX//2fFTdGeV76f
vhsHm0x8SgAgeLoRp/P9wLAF7DpH5USZ5aRbUxYEFAxLzJlSLn5sPLgzNuaS4ihN6DAt+4YNihR8
aXlEIVp5uE0beczp0OmXcGlajgjwDdsFj5WKwTocjMZ6EncEo66ezJT/yCw//1oIbRdsczJi3lJW
JtiiZJqb+VWSBULLgGOSTPvWF+W+naeKi3LauHmBt3reeM3V/51QRKvm4Mr03nNlvb3Fi8DJwCQv
lj1Cxw90mzWNqY2f36cZMavajMNdOAQRcVKaIwVqV5XiJ3FoyCLrCrwzzPFJPxId3zIAHeYm+8p5
eNKfIopZOOpbOHSO4TuyUSoADYj77GNzf2N7rEXLbHTplUt7BugCjXUFU++0YOZSDhqQx196b4M3
Nyo7bCCp6pKG57D4zGrx1LjFWk6eB2/mMestqdu06Sjv0n7y42LPZSQ7qkc06awFySFubPHPO1eW
jAi6GbFxxN/YT3qwjH3uaFM1LvzUcoWUL74qe/w/CLs0xC3skh29m3gywoxXjbepjF/mJH3uaO5r
iRXa8QVUuPw2vWYjd3fNC2lUEQEgULSe8qAQn0VoHuUhELieR5r++lUCR9dewt+x2kV7b3Er32Tj
w+zaGBGx40Vtae3EEyDs7lYx++My/bMS9sNGGm2pTcX64Pb6FLUt1D586+A3iipSroBZxJwINxvI
EVbQObX+bZQ9L0b7v/v3h4KUWsmA3yFM62QB5UbRrN5Ag/BuXto1d/SVll/fg9tnFLKos4ADH4Mv
Yj2vnpU7MtEAyVHxYSjmHJI+XvIblWJCRqKywct0VoNefgNX+59Qi8R206V5V+B2DInGy1uTlDzl
6GcUvYsvpm3msiJ0YJvtyl4+ur8543VS0ePhniF5PBeiqqB3xJRWRDl8Gk/iBD+1mRHkXqiL88+e
TzddA2L37lHYAJUR1zosbDYtmXD7PDS6UJii33zHr0KxlOi06oqBfToPR+kOCo4aNYidfayiMRdK
a3650P8oKiSu6pk2m3ZLuCuzNIfNnWQEe4Tz44YcTkdkK5NfQ22+USw761F8pkhwpTl42II21xrr
HEKKY39F3QaR2Cynfv6A8WTuQZ2vqQlT1K3eGYcKWKor4NB4lWrRbEAPkDktNfrAF0bhYQ8rntus
lxwoF0xHJhvXH/lRrhMeVWK2onXw3ICcI0WWeI4SEf0BSWYfFgaxAqnrBISQlS/DQZbmBK8NFcZI
mMXQmdkS/OfOAy4PB8OaDuWy8F70qIem/KpNnNXcvgDb+1OWWGeQtyt/juv2GECZj3bVjliYyq3h
Fa5XM63T715KuJJabJCViHQ2Z1k1Sd8CaQ80cMFf7iABDsWBcVkEA9YxGqCMvS2KEyAPE98PQ7/C
D7tZkWhDdT/D3TQwYcPq6rJbsfn9seRRzw38iIjxUJVFNsksfACKWFyRaxIqSWeqamX7xKmDNo0I
S9MnFWGHGDdPxhDVHjdLVxzJCvsCvumKLLA41TN7xFy3NAWZgVblwr9cGGeEjL0fPUMgDKzJNNmN
7OpGz3Lwi3A1WHC1fO6+lY3ARbODrfDkZfqvZLDCJX4Xxxb5oacB1xYYvHZN9suXGJ7vIHAzSa/F
FxQG9OkpsvpPdqBAgC1ERAAli0MEZbDBXTHZXKWgMsFYp0CIK5JNf7YKmtxzn9luZ76l6Mi6kVgw
xpuVC/6CHdVHcYmCkVM6Cbs/fCUR/s6gpMkk45asfspkkU6lCopOgD1G4WCvKnaYAPa4Bn/XQifA
ShMmDBvH2CiwgwNzOcpAPQmEL+Fn8uiCF1ZtctzCEXOjI0+r6hVQ55Gy3NK3MAr4+G933PaG6J/M
rryKNA+PfJyWLTIqYDlyp7f9CuG/SASz7OwD0c74bsaM38hjzBH+q+NNafsju+CKtkAuStZg202G
cGPn4FiaIp96v/kXCWxWrT/BUHhttqTDl+w2npEXG/+QjNRS7T+7phjpHV2poKjl4ZYiVg/0I9ss
80Al/KBzHpcZCvWWbnHvtKFwmMezPj7MjRSZTZKjGlCTxRdnv0L62B7bDOAo3KPHpcmACsIMhAmH
Trcea99uwWs01GUpcjCtATXKgHWi4oFet4HXloa6LcXVGelX7rxusMlAyE9Jn/zRlfvLgua2L8tB
R3GG0MpUnwZjHE1VqLiPznFntEfMCZiTBjfFoexxi+th5+cE5fuVgKm/t4SAhrTkbGbAUKFzvRQt
bVUALya4nfeqzo7xu8c9FKhWE1l5m/aRUZUx28sugExcfMPRZohcTLH7vjis7kpjBTJIHykHF68J
fvK5yVokBtyCp3U4/pTXckupigu+pLZsncY+lTR4RHJDXqcHPQEGC1W3R0Pfiaebd1QaWCMQSxHV
kjmAT4rafimROs3Jkf15G9kisTqKS5V6HzxypvlJcvpZeOLnyHCdCiuxXXiRDJzv+uD5S/G2MovO
UsjtCZMtrAyrT4BRXzsTAfjGVGDtcwdtWLxBf410vGVo4Vq/po5yDGmPYt4xRHhqt/DjmybJOT13
g40tFku84+5MQPMg3fydzXMngRe/Gau6QM+U8EnXDxLT7RX7tKMdXLbhTth1S3B50aMEXKrxNgu+
Lo+6QkTeQaQVJq54f0/6VekQMpjHVoj/G+9orMcTKV4WiLLeMAQdTXDzo0cBwVBxDvKRuvekXkl5
VQovb7R0ve0Ayr8ajbeXGL7AJoAVRAeHlPfW8BZSW6PQBdTO8e5cKlx1sP9GlQhx9koOvjmU10hz
Fts4XNui3uZVTbrOH223hI9mbYFPWHTHEKU6Cb9k/KPdMCMlOkLiY++S9zHEIDU0ikDsaq2OPptt
UJ8JmeyVkiAOTb8/d9URHzaD1iImjgVsgVHr4iCrZBU+GDPavQmaUPB3ZX9t0It0R5zRYfp00Qk5
CGfDKvkcmwkrkbax+cz2xN/ac1Rme8M6paqkzzyii2HxXDUTkPiJujCxUN7u8vQFH8U9ZSFMQGQG
CHjgevrPml6EfHbe0MjsvZXFkJie7ZAxIx7s/TNNoO8FE9ivDcFFWwwK/22issDmPWEPKj80Qtd7
p0lzSYF/k5bmQTblytgMHnM3qTZxBNj2PD3mzH4/vTApuVW1E1XUEgKgv8f9btxUkS/7lfQLcDbg
MqD3AjRmaYuG4pDPSyUPQuRI98E4X0t2NwDvOI0t36SWrEcvCkgrdqCG8R3DJNmviTa1gKt756Id
nkhLf62MdZEgJbbtuZy6MZa7Dk4xYEb3wRD4b2waZlQwzcOwoU9B+wXHBZqFboas6YdYv/wy7hl0
K4zP/+COl1XliwLFiZiq1iUOBwXQkl4o//hHjMJkLgufmc9FwdxNY5/pZ4TKq21Ai02j8c5FUP4W
YoC0KyjpgMxIMFIiquM+b39ZBszmfukS5K4VKzpaNj828oY7sgd6mo5Mb/7yHgPfqTntZOGDvyTm
Iv9LVTPcoW0McU53w2qvDFdZToBlHreqSp9DLY82+p4Rpp+SqqAzE+pI+F98+a8oqBfSsvJoRgbv
im4Tw6DfKF87KSAvpT6KsK/ozKFNQtXUlLeiMK2qSVEXsfF6Y5MqHVhxJRvLdwC+OR2bXdCTM84U
HjgCezK70AM8i6k1EqfXppVHmBaZ9ETHE/jIgK1ZlZQODWzJgF1InITS/gg9lJ9ya7zMO/D9Xq2m
iAg0Nz9XSCGiFg63ZzV1Rv/ih0RJoUufP9CS2CqaAMxYqmjepsEN8ZgF892kjQfRKMCevA+TC50r
zzgHAEdrNO3PATRBjEwbUEShEHvPROQ3d1zkSkeXyMlo05M0JmyQo6MSl6zeDmDYtQMepZ2LcvRa
sp9ZUYcH7miJZYqCckkf8KnoYaDAijmKRsEM8QIizPsHofuYcVI3pGpEGZ7qeVBTdgS3Zge/OANW
HVAoEjRvx9dEVxOcO6GVztilYN+YfOYZ9OOYBwTuOkBaBTzacctUbJzYoTrIdOhxImmUAzR0XZ5q
1TxjDh1tWFeZ6EAsZOzWOjJ2Agn832Kzdnz7xbw3Tl2jEYNwjI5z8r5JXqIpkWvQf7jFEsKX9L+l
IWASzk/izjNi8mdb33pctR7OmG5TNOrGtJ2FEINFFNwuDzHI6jKCMxBQWScsxXmb3cz3Yndiw4Eu
hX/q2iigO8DDW2Hx/tpzS/VlwNyoe0u6aqNwSkI2/7wqTiPGSSIBRYwGiN0wyJ7xi2WrTC47rGFK
2cjRRfDdNmd5//7pm4HIommJyure1VYVt8MC7n5I4VN66qASWJZS2ZjW1RSQfJmKZSZUcqKEFrCU
FZ9LKi9yEH55aAqxOnsOqWR8F9ZCmJad2hDCv3UeTnsg1bNV6urHH9fO9UsxvvtQAut3NuX5oxx+
N+muaHyPOgtF9ulrK1TiCRqVsezoIEsqRGYwnIbTrIjqanMckDaS1dTbbST0289L65xKBGzJShfn
GkBbuAp6sWry/JBSao8HfW6RpxRBRydweyLczaowPAREFVFCcPsyU/yO8KQGIEitI0/M/Iw3fZHC
7TRUAZ2VzkFNUc3bzcSIQv3BdqMTZz2Yfl4GBvgPB31wWglNm6Q55qJphPDfSysaqFgFzq4jIZfM
1ZZt1aqbesBeXG+auDqegzoivLbbgHfd27gzjBqxUfR9PRztBN3XD2OvGseM5fk2oC7ar3NroHu5
dRCAFd1WBhXYrzdsahs7C9/XQQKFQI9Ta27pnlgMkU3PL05jHo4iavv7aah9m9/vEG8Q82tbw447
vlmGqyiN75RYzoLMqCZaRTOfZ+UP6Yu/5rcWggo8Z2z0D/S6yYVUse0dckgeBX40/JfhkAeZVy8B
ccsW5GNyOnqM4DXFuHvxA9k60g8KgQwuPPA4LfMfAgafa/zcb0xVbscc8I4VePLmOgcQNN4ZhTuB
RoMb6I1WMqM93XZPq1jS0iJgj9b3HPg/uLmhUVNlq0UTwWD47FJxtkRrzVLllkuMNcaaZOOQC901
lk5KmjJtXtdHZ2mtchrwdl43uiAB3bnscPsm/t77pJaObNsEXdz9xGEMDYzilFTl9s9vwp9fz5LJ
89SbnLOxeZIZaIeNToNQ85//DhZaKgw+/Ed1Ze48pOl+UQfSfnB7fViV6RMDYHNtuI/etDXqkmNg
gjEufVEavWLWi5O1cvknWrV9bMvrz8D7uNV3Rs7rHj8ykzrMpNmGYh235N8bG1KkVFeQtZ7y1m51
e+UMd/rUbTQSgrSA8ERb15VOuw9wjZ6InS/EuDQiHTqUSooHEPTKhhGEZixcL2pqSWXxver4rSko
pGihgBf869K+gjCtcfksbijYsuWNVsNeNd2kOxnJhrNDys0eudW80L/PxPubFfoZObL5fBW9PfLs
0U0oPk5ox0vR4nm8AmOO7ipUcOt7REIVUNPx6zN+2S1amsiDVcdvUQMn/ReCf7F2L6bQRqBJi0Bb
FTAkvm5F/CN410yKiouR97KMNFffAEMs123zMhzpetuyKIDZ2c2x3/PcyCcCHL+nN67NKlVQcYeD
kXwBWd12dldQ+QSp1nWvQpyhli2JfnTWIAhsOS5QVBiOIZ3bLFbD8NGur16/SAeEJpc+VO/4Xlhh
+XWuU6WCxiYzKvRRhJSU8zdpPimzhKdExMGQOv+QDNKLeXPIzS6h0ZbdRuKhhNrzrhpi7IAySTFa
Pw4OKIhXMibZ+wV6d3Khx5hZcSzsjbPIt3SfVSpKJ2N5j+6dF+BlKvXYx2R9iM69U8zm5LagAvcJ
GfpyoNFFaGnzjbmzf8Sfo1N8+l65EnGNQf04yN4i2HjcSXy3rT3cI9Im5DdWJxOey/0yL2pMPioM
NlwXhje6p/PDFlP9FKWbQwo9yHBlGrhOzXRiCoeITEt4vQBPDUXJfMeG2b0JrYL9e5ejtGKd0ndS
r1bMifIJR8CTv4g4IEfRAYjKV3j8jUdq4BZUjAy9p479WW6obT7rsI9YAwJEO1pkZZlW+DpAUrDx
sZaYF6Gcq+NhP8BlKHbyoZTFWtxS9bEuycm/cpCwgXrO/QNKoutCWahO4QKSpsArnkXYMjfj8qFF
hyyz27dIpCYQ+85ZxfwwO1ryp14mW2AAjC0QmcWQkWJq9C9GTQkGfmYMcdQDrQDIbxe5IMY1uMdB
RIyGQQdII+ioTxzOFqc/htt+dU3cgWRT21g0Eg2s6mZEH5U1Cvs2haZrHTq7hbAwAdA8/enBH1Wd
rzXBFtF7c0tGR16JNhi0nHm6R3BPPyugFdouA0mhTKmlbfE1xGD59G6s7tJWGUsY85yRXWDr8AHv
X86CLnIY1VF2sFj1pJSGO/mJB6ACx6Llq+g5bwJkV1p442vMuPaCbspA8Tth/kx7kz/e7S3ltMfA
HcBrUz1p1C2n9vvOKCd+eZv+1qGLihU0ABEUvHAqzLymlpLZlB3Igx7oP5KoX4zKVHUejKx/Uwft
hF+6gSGh/LgoWwuin6IlG0fj7Kqzre+mxOs+y6N9ryTnZZAVeMDwxdRlyjEPnNy6kLNDTMEAhrU1
0N44jyBOU3/rOijUI6FBPQzuzK63/LoyesO3qGPdnlPMmhNGb9CF2AtcnXl6eRokWeqcXXadJTbM
YUof+zppQZyuH4RAHNU6QF3VNFL4n4+D/9/Pr8kE+3D6P1PVTKDdRLogJdmtktFeNmrJ5ufv3iZx
pnSQeYRNkWvV0fs4185BRaYggAnaSJDVlHI7enfM0+vx1U7w4l/Kdip4sBwmZC34LaGs2ma936Mp
rxRcQwFW4B6nE8/mOm8IkjlFLOCIz8veV0YCG5x2pTczZw+fP7Q626e7BpnwQooMxCu4/hpqi8zm
arJNl0o8/7imx14xp3+CR3Wf0wZR118bIX9yfm+fKIIIVllWeABbf0ODYZpEcLLfaBRSXtpWDOtY
6UlUaV2DswT3uHOudNGK8zvPYIfDd16HrEKCw+lJX7jgqnZMCjgMeAa8cKrIMXhUSE2sftkreF34
uCitaXMzo5d+h8eViCUvriwqRMeQrqZ6UYnJ3eyOJQLzSbqL0QUko7fj2hVjEoO5BUuRU039kKb2
ziCRAqRyNkGSoOIqSMdQkg9J9vSFXDLxOWup3wDLxSDXr8v0tXHudF4ktMkJOsTKJl0/xhpAQh+5
HcDG7oE88kZ3sa3MjSDWmrxCim5hFQr+bxVVlPUoalupl3oX9oVPas+ym7pEJ8IVJOn7hMZV2c17
pQxEc55kC2cLzPw8Dex8krMEAzLQ2YqKXMD0GIfmKHOYyOpyJrRNfEuhjKmVtqEYDAm+u1/DVeNT
EShguTxs61lSJjs7hFR8PsMu/d9F13O2zfKpStPKn09PY3fvDr1sDpy99ajIRoLEsusfnmB4hBAR
S2fG4fUMdiAA30mwb3ybxuAIaYCvetPFhJKSNKqv81IlyMaFYnjldCtg+MXTxs4T5N9P54hyJTer
GfW3pf0xcVkVJFHuoxL1sClW4905in4qLEZv988tuVEGigSdDRpSAS+ha1dGx+gxpW+/raY/moOc
k98TDegIb2JnxGs4WJw5PKr8AU4mjj/Rvu+Rw8MEdMvD01zNEg7TkJD+DFL8DPN8wPJsGPSBg2oV
+Izm+IVCpw7VMbKzWKRCVdMyDn0oRGXfMKKfsudRxSOlQzHki4yupZYTfizxI97OHRhRe7hqkgiE
sPstzbfjFznqQ97WezaNmMlH582ONxIyXPXZ+FcGnCZgfOadoFWwyimM304hRd3XQnz5SUKTgP0S
zphTbrAwnkJ2q3j/oAl1l9omgGYtKoejuqWqJzkv66GX27sPOU97APE2nFxXIiJz5pmJKkDjV2U6
ucYS57gwdNuI9IaCmMnCJSCanbM/+xnXe2fpBF2rKoTNJkCasU2q6ErDKKcgRuuCFBZcpPNrxsOT
at5o8a2WZMeczWK2rJMJshCUka+5BN8cF7sI1ncEg3jkIwLAJqYaPDQrvxckB+SRjxmAMR0u1WlP
c1O21Sv0Bp2ru8GW2XjEIzOTrS1jiPw2Yj8OO+g7E5TsrAH/MzGPgRpqz5/BMMziBZ9St58SE1gy
BACMuD4ZFkHkA2Y4HV2NNpuccHgak+ZKf0YR9MK/CX0iS8OnAriTZDe2hSPKlZmkysngxFH9FKVW
SN0Dmwg2BfmdBD0xmnjXubDtwo/MWEBwZ0gXU+8PNCvZJLTI5EvFTbQvlsQBXhMvUBHVAmBfs0Pp
M/RrNRbj4j6oN3SwvScIMAOnTv34dDbaAmYgaijr7OBRbiBeos0fyU1L1OqkoNc/GtBmw6qXRrwl
BFnGORrah5M09VCv7/9yVlsu4EARv/30OrgdfgIKQ8NZVQzt1+s1jZOlgscZk1yBRzVCN6jIHdMY
+a/xiAoiB0sKK3ar+zBnH4L/9B8hKW15R0sVdQojyNf+/H41h9VysNDVQVNuQ8RmP9nt5AlwMBw3
ASPmTQxtl4lLnWKvCV2mAjX7KqnZZw34m/zidvQNixamE0p/4vjyx4BP+PufbndlBMxIU8s8Ngju
2uzl7fYs/S2FtgVHcYghf5XXT29gUyQdFE7uZziMO/SllfU/9oOM2vRd8h0SGkCEgg7Dum1wu4nZ
PDF8nPPbTNuUbKG5PvnuC41dHiZ2didvrPJa80m2eqo12BCNgvwONW+t74cPXqmnE05HThG/30sB
eFKLqtT/Q0rggjbCgVlFjuGvfv09MHZqIA25JeecdkQiy6bSakqXwCempHHGncQJnQ81QDtTVmnW
CSWnYVbG8ZQ1usXQfYDeFXzURcPC6YEQUsZI2AyNVLPPJMi89LEpAFYY8eQZ7ZXN5QHqHZhTevpc
9VNJdmprw2V1cdx5WY3AIWvRCuxkZqgu7xUDJJfC5CwJTfM018ex4votsFP9l3d1zmoEq/FTrkoV
yDxSXIpqPzQOA/oQmIPfLE3IlZINNlrcT+mXMwLonJwE9CHU/9gETLZW8t09l9RbugNbI1ePA6GU
tLnkLOfFMOoKi4L+duVmjvSnjqA79ffmEOPd5h3GEb3YInZRDIqHrVltgUeU9xlHxYue5j2jbNi6
y0Pnrh7RTGyE+zVqaZHI0L3czsPdnS0df82L3NaY+VvQ50Hcd32jOxV0AS+R3LxADcZREKcLDkkP
RR3YGj/6i5hhw9gfv8SVQs+oHE4P0kSxTwx78YoTARZ8HZzRNg1+SNEf3Z1hE5sudA/qTbBpTgq3
mTXjDpl/qI9sC3ezUiQP0vlittMu5pTNPVcGEolxcI8qSJ2L647aiCntSrK//7rnEMmrPS2Qlgk7
ieYS8N1/J0OD1lbUwBOBPi8POWm2CdEVf6C1xsrldvYzz5MmTESku/MPZ5EYGVQR5r2xEeIgSRFy
lXFeUod2h3WpEzBUCxOPHKnH4nDNpHf7/7Gm9fLAPIER2+DvYkwaNz1DiFs0qFdtvCBhc+ZLl1m4
IOPyYjxe6S5wehzek/qKuZNnR/CTR4S1o8MbFBk9pjHeCfm2t92kXpUuRiS1N5gMFwU1SOwZk5NZ
kUbZjBEIzwDpcoprslJ1ntU6xSx24Xmnl2IoBjLMl4O1di+7/WPRzuojdiEoYnTG9jO1q57/l2k/
eKbSG+2BYWpsiWH2sK2nfIZqtyAGRZq07byxBQr6RsRPkqvzrCjj3mMQgnpIKHM4xJWyiI5akIsS
H/KErKdx1pxABKeqb76tCA3loDM2WFQgjw+pOabq199ei3d95ugCWpF+P5IuQWuGL5SS54AnlYuj
QK8M0pUEpz3ryzyerFfyyTG+qRj2YsiJJ9AhXGFQRPht6UULkBdF2jqZR8+MpRgyqF/wu9qvaE64
xIouxu1OonbX8hOrx7w9OxkmvDUVfujb30lNeryFROH7Yx1laOSYXVp2B1v0MSPkzX9KRVsgbx+b
v/FtwhxpUtqYENij+ihJOHlLGniHak9zhiTmfIA2om9Ynp/B2woRyoOLvF8sRXAmY/wtgkUng99W
Fjuj+n+aDEOuRN6vV9euFVa7SWgqA4LKJQ4bawl1VWqtPwV6VUZEpFNopkORYj+YknAecE+a0ZEx
akMPLPA/4xwcMYbevR4Aa8MbponciyzLCsi79kAPQw5YPEebafrMi8jxiVjEBpLLjwIaSkJT1WZZ
Ubw4p4PMOiJgK2OZ5ephhlMBllcXlWoD6Roc/PDG+O3bhEFOI01n5r5WXTpbMLmj/ixmFNv4tDxX
GG6750DvmgwndFz0vZjrtdVUJjMDJtdx3D+odnClXoFXiwBDrMY8SlyJa7LVuS2SYrfVfDXVrwak
BxXAEZN2xJFLQaT+odeP9/VkQ8cfnZvE2zdTp3wBsQ02RPkZv13AJpZs5jzICDOQJuC53E8/eki4
zcW1+7Wo5hpZUYKcd/YGuAge3WLKc89Imox0qjTfOi4/k/lHg2HHeoe5qDrqJCLQxkyqbi8otQMU
OyJMZPd4M7KfCioldg9DU2fbjTlh962AqMSmETONc1P/YVbzcGP4uvVnurqxW7EqZJIj8CMccO2g
KX+GC8aDSCcBjT4+2ECmBsuJGMA9x91VQjqI8o6dpkvU8CXmugrvTOt04o6jPg9Nujx/EwWU/rVd
WYnGjayxJ4+daeCT8pDJymGL+sJHG2JPPiPcbtxHguuKrq9uJWJfynxagN5G47AtlmlqBuU+AE43
rURA+NhIxfFCwRysCN2V2W39BkIhHt/kiXGq8FqyKMrkvdiK9BCEtFJoXbJO8B70Rl+ZEsylbP3y
IsfbyqK89zJDbPQ541nJVQCkEeMV3Tq5n0UMJz2uSsP/Ef6TKEKDtIqd+ntEZb+WxMbPfygcG7rb
bJne7fl5Q/naD3I3+5mEwal7xOXJ3XSt51rrJPLb4uhsRKPlmMAWjjcIDw57fvGDOOOR+fkcqAcX
252YqaYb+ObPL3viflu1G4GgP3n7CBOiNUNcnQFnce1ISZTkjcJd0oL0cXVO1WMGAjK+ANPPSzTz
HHKKt7vG1bJxR1iDGouwxwa4EPY2m9ai1o0Aqd8t8ZqlPXq+ABcS9OqWLVG0kQpB5Rx324PhtPd6
Fe6EmM3SC5ZmhpraBHB/c9uYb5qs1hP+X2FFomdQ3gVnO+JbNeSB8yST3u0zOOyEW3vmBqT6TIv7
byVbZHm30HetPh1wfOczqmKTxZ8ztF8MXSF3GI/xe3NS+R6QNyyYx7Ddp+EtwjB+1pyM6g3KlEmH
8+gZUqWnSNIJ0fSrWD0dveUDErJcjPkFGRu8sFZC/ytrYH6v3EUcwKII/slWaj7bGI2Jsb9uxF5+
zsgQIDJ6KGs6wVBHol+Xw906UtrmSie1F5d6xUANsQNge2WpFz1RHgfjfU2qnIOZrcuphPTw0JG9
CW1Q5XQhuGLPhO+RXLC7zFSwGSDPchstlZcKN+fJiGPSubIDcOIFmflqQmKbhlDoqcKgxXP52l9N
lHXAbrku22v3nNDnAXhdmCj2hgd0bl8Es3r2y1j7n4D0oXj9O3wizWYNelnQTWzXliOwknelFIN9
2jyaXvvpIsVxU0PdlhrLEwK7pgS69Ktp3y8KSzuBNRha7FvKK2I4GO2MTg1diu3cODhN2mX9ayAr
s6oJ7OPS9Q3iEBgDfJUFOU6TT53AYB0gEmQjXVFSaCihC+XJcU4IfowPr6PlMnFprEUBgajVu8wg
Vbmc50Dm8U1ZsKMH2lEgwr1qZI/ioHdNpG0cypUIrGeIRCr4tWLhJ8/OAApmYrppfuRTFcBRPIb9
3bIJFhIg+qF3R3XmaMlPJUDn7XMJpuAMp/UhG47S+El/xo2VRInMMRlPPp1dIHw3a5Sa3rv/7y36
tG4+8aez7h5kGuf3mMSzB0BttSp2hwxW8xLnz91DY43bSuo/uXrWVHLKO+x7PH5ZACCowU9TtbFm
BmNeQtVxqyZCtlV7EYAOFZjLMynaKL78HOxz2zWk7MbTvvZ3sJqtBV2hG0X92IgJplhH6061BB+y
n5QJESxhJ5k0HtID5F+cC1UyatAAhK3Jqz5pXm2uM29u3ewzuZjo6iJlYbbPg2DjS+Ql+815zI5l
/mFqZn9i+dGBcnhOb+MYr/WciCIcLV1T/YyTGhTmQzAy8QqjQbQrDmSJbI1uWq5qlmBwo+udQfUj
VZZNfmOiiT/SZG/miO0QtNRpsFWGSb61jlIj9gsT/Sw4wVa4SSt/YMHctrlJFYxYRdLdDiB4DHbN
iplBf3Lhurkvt0M27pYjIDQqPKTaRG/7nJDg+T9uCpYTs/Rv/4yJArxQ5e9KzjpPxqpQ27E2bXnB
4zIupKEkzfaZkH/Du3PoHlEDHhNKz9jawDwF74Z4o78OmvqeLLgJvTpQO7VVaFk5lnFVaXKyi3+l
dRYmEe1M/5Onq0uFs4QIfiWY5qdbIv1/cOJmDJYiJY8lib2sGtXeg6RX3WBnHNgn0a5IV3Amz/HJ
i1cujnLKitzOsK2gi6P5ocg3+I2RjVY6X+iLiKRk6ZOGFAbvujPWb/d3fiSPnWKDeOVu0F1Gxhx9
vurBYaWMKk1G+qeaX7y2/s5JUXPvD7IXIPSK93XLHbMHjMKjiwLW2D0oVdryODdoph/16D7MjNJW
s4suExqK7+qNLB5V1XzkHgr930ocOn4U+afTQSmJRgqhQoMwaqslFkCNMenW1bJ5csCOk6movZib
tZzJB2nZ2oMFaq1o8tni7ciSZCBse6HE6mdMWV+MR2Lt9mC2oOsqcBqvYs1w5WESLFKBveveYxoo
NjGvI+24880vJ51xGtU0XGRPWzN6TntOXWwmMMydRinkMkRZUZktSB5flcmfbQVpClAfLrAMaHm/
3H4hmRPiLfLxhgBBu/JqmMdlLdTKLdNa8nZSQ1PWqc5t5v8DLijaqnygCSlNKC1NbUT/LpFNtqhW
Watm2UVGmcyUh/W/mRaJrGdWA15LcR+wV8uMPi0KbLXeHgeANC2xDgMUQMJwo3eoTLNhUtQrLfC4
n0Pz43DZ9cDqxGf3E2FM4GIN4zGpXNKyVT2reriTsd0kG5GRwbFI5/0c71gectDTMsDzhc0ipyMk
0oLpoxn2BIxTaA2hnZ/7JpmcJvWIN23ir2CzOmFI9Y3AXxI0ZeJORu0gxDV/myYh6kLdKYYMpwsG
fh2zQska5sZZ3N63I2ciFatFj5Ce2bkhOCNF0uQP9edgisgdBHwLP78hknnMvqE+yeC78MZExQPG
D8S/hnZJYPVNjDVkd3k4jLjOuAqfvpp32hhRmSCSQz4YMjGn9OhBEy1tSo4WTSZotrDJQ//c52CQ
tTyOZqgo+Cdterbvls/kJK+fJjvQ+7IRuGEiJ6ijcA+zWy3NQVfHfIk1cD7e6NHE3SrnI87piQM2
kIwi+QarO7+C9+5BIB60dC2IbGX3qM1mttt0D3KzA4t5hc+zpI6cFB5FhdU/s1cebWhYnkD4NtUF
ZiDTRglNO3e+7KgbWKUAC2FBq6PU0CeUglCyErmOimVSv7LQlH7X4d3f9KKIQsS2M3ySE4XAhwhJ
rrIHKJb9RY60TX5I29KYS15ESakQe+J26O06x9XQcfnHimtpvdOVkWFXEeeFvSBiFxXc8pWo/wo5
oHErzjo+zviPH9+MDtEl9Y0tIlV1KNTQ5ITT+np9oeOZPexFfYWTuDIkJR5WalkPEV+XfH6Yv0QC
blj2dRADAlp6D5+ShH1Ca5NyzUHCKDYzHGzb8/iLgE1TzXkUA1Jq3rhuOhE3fGFLo1uAIDFcIzB4
N7G1PNpDzlxmHm0wU/FkAvrCbXxE7mmtkWCQlAnzybBjt9v8UYSH5R0dJkKO7R168IEw+Qx2rMAG
yiM8uDbJQs8b+JUFtHrVuQVNysIxZg5E+GKAC/lj88rD7tffnJhvwuQxJJa4EFeUdO/WdQ3Azm5g
3Hh/wu9WFckM1Hmt6Ge5kF1/itXmLuJLDLs79uK1qUiigsWzX9b0SKHCIuQPcSswR5nn6hu5tbDU
9SLySPacx3F4OiemzoX32LART3z6bHNlGnV5KvgmYZUbi73SEb2pJBjRlkIADwBa93HkQcev2keb
ROQYIX/oQy92FLuIDre0Mikxf2i62zDEfncCersJqUuehdTY8CmZo3UFfJWM2wCrLivRdGPxI8yh
TRP+zW42Yke3jZKMqUwJSM6Bs2VPpMDWHoNhh385AGbOXkNLJhJx4hAifEd1Cl0HlkMHsW+LEOJI
se08X/J/vRDMQ+/cUOwvvrd5+YmA+wVkr06X/eAJQ+djdy1XejPAdTzGSxGXdLWftEh5Ae9j4rx0
rTzMGKNhK0YUTvwFFa5+kIaStdZO7Gj7ofmVS3w/xZbDDWks+LthLyHneuxZ+m4SphqPiUCVKDRQ
48w9g763MWHQnD5rH0k5hvu0wflS5BSS0SMbcUn6zvqf0bAH4IHfiMDfCFEZaoWFIy4Hd7Frf58K
QZh/PQGfZOxaaTDVrKeizb+OQLUn7JZGjQYSqhqHx5Gz7fjRAHizpxtpqDxSgW7IT1ceiMz5E0gs
Q1/0CpNxzsin3SwTkK/ZcLqTn0gR9YFWfU4or8RbYA6fWEqsA7CdZKDh8a6lIG34lT5piUicivU+
JmHBHoSeNR/QjvPLrjE0OCiXy8WZ/URXMCIW0o51zn5WbhfqjLe96PdB5fLzLjYNDDZ1owLKAU9m
36cJIfBkZNlK5CSQOals3BXnsKVN9ZhTBYOo21e3xxi5g8vWYWD6TEAoZZfNnxYleA1LYlaY1Vw1
H3o0krhTNw296Y0Qgx1XF4KnYn+AbhHkqS33nhXT15DKp2GgyWUCzheEMLyVhClIBZdEUvFRZQeK
wvvfXGco8toB5hX+qeaYoubRPaJD+yS4QFq54cAVsNnbUqC5l1aem9k00H1y2/9VscsnJe3lCg7x
oCVX8xXrm7Lu1+RaqDZuFdiOMEfskmGNnUPPtvaYvWg6uSS3NJy1vEAOGvMvjjemHH6pQ72DiLpF
ZLEJIzk8NOMsEF8vT3OxRgDo6iBJ+zGh52kCAcp/2Upa6rfoFaK+SeO3ARgnUSCZvADBpF8wCDGb
TVOnFgRiAsl6fj71UIh4cUjEGWyOo5Q+j0NR8GMgQ/MaHmB85bRmPistTQ8PToeBXnGG/1EsuTqg
N81HPOLl2UD4oYPhKyBE4EXDMGCKFgd5aAzKOCrx0nST+nzR2xXHpjmwHeR0efSQJJIDQm+A6ehD
J4ZmQBmSRXA6Bg4VCUVwbeJYe76gxih343752QgCFs6KBFN7GraUcKZb256PTzgizdie8B3D35NF
j0t8nS+P4j1ucZGC32ZV4hKD3EC35RIYw047yIDvESC744aeB1sgeB8APVtcX0WyCO9AFvF7eHEn
z7jMYu5lQJ+v+RcN3zihNvLUoyupQkRpqrhwekZHv/qldQtmsQmaXkCYOWgIFMRsXpONkiwtWC0p
UPm6BI3Qsvxl6GYZXCFvj/1QRi7OxlgSTEsY/PgDZuZJwD4aexciWGSU6hMAdlr4IkpLDvcHSiZO
DvmOgDi/rHyEa/ZK+w1bWMnTEEzU9ijpcPZdtROUCyV9wjsKGT5V3QVH4R/dS/QSRxwUY2cBkj+Z
G0haer+ttvQg+59OpdEYgbS9zoaQK9OR+qSNjmKMA8nOj+ZuUy3leg8D1/A6wkobCyb0zmW6CP5l
X2cf5OAygJNGT06jK5Lzq4Kd2b7VRSjUmFhKeGLoZigU1Qu8LQs0YTxATmt2KRj1xjMo1KfzOIvf
QT0lrUyjeBVLfhR9ikbidEXdi7yQNteuboOztiARbevPoZzpY1f+dMcBf9NDMt867Y9WJPvAe5OB
olgRuvuAXWYBdT07hSOV5U70Z2CzA3M03qn7f/Sug3JCxfFUO2AznCVMMM/6hamY899i4U3QnMXo
Jnz+W1Y6dbYH0vVCCJkUCey2ed7dLgqnxaqiR1dV4Fj30xcC76JI4d03gDEeH7GtEUiUOhRlYGI3
jhRwZJahK+q/aavCZaRhDOrRIYtqXE5iytMVtEUnoEywKJ6wozHSFXfTv09xxU/Wq0epa5r5gQKy
Qo2Xl8KPlj0z6ILrbr/w0DGcIie3c/EqV0VBQmOTgWIWud8D0G+WCEcSy8YZ1eOI7YsibSoiVwkG
Ii5BEI0mo5D6W3PsCMtxnFG/pV7nucjeSehNZsWQVdfki6C0rYGwr9AKvNRZSyUWfr7W4VVAqlOI
210vEZ4rbiuiouZN+u05L1AOUNrXZ6VrzJ2tXxqmgBoMUtfLoni5KPpu0TWlk/GC5QNYpFqFAZlk
Z+WBaXt0MJtgfReBHGjfiRqU8zjLijxeMAk2B8sW9389FiRiMNnctD7WbhVzpPtWIr0yI3idKXFw
SMZyAv46hJGUb32NaHPKdwjOFZhFKjLVzpOwCjsXPc1YMpJoAibxIPGIPFBrSoELXBd0QdwFXkue
SRfq7cpaoIPCz+Kc+CjDSyT7SbU/0CXmGSj39kskWDbHhdrVY1legvkdQcfN36kKPdUXcwFDFjV5
gM/Gt+NpezgKtyq1c3eXIqMw92qS5FGevn8GU3+vQg0DqsVTLfKhgsefCVXjIKb8KuA99rGPDBt7
uwvrsIpxY8q5geMWtGxOsIsPbOteApXaIZ9GrEsVJhlrE/1ZnFaX8FyZLewix7GY+W1PFfkGLFcI
7fu2Q4KewBGRIOBykfxFpkhkiVcPWynZ7OZKICmZ80k5KEVziBKTinoczViyDZ1zMd9A3+AouO9P
9iPtiMKlor3uRRjjWiMahg2smE4gWcp+PznNO1ugFDKnADbTkU41+mYGXIZaD29QcAo6iTN6GA5S
wUjifQSYpQ6yQDmOohcatEGmvp70eQMSL/X7uwtiklqQUn81gkkinL5iV0oAwlytsG3UbIzHc4NU
sMT8l6SOvd2OyIvuCCQsLQkjdloJJepd2weutMEr+sJz/t9v9nz0oTI9v7Iivj9khnUd/KdEdG8v
MnhxeWhP8/yAahoVszsulNtDRBLK8lXua3PGZQdJ16XJAyPe2rV/J/gvx0rfb49Vl7U7YJlpsBlz
ykAWdxsQYlTq3ElcdyCQlDp1+e5qpD2CM6ZC6vqmBVQ5KOjNKsoxZ+/S/+1Kmg5dqVV5TXb1i0ic
CCVvz9FMHPEKVTen2viAxk/gmzm/lQ3nw7wO+q0aLqoiGlFuNHda7Ki2kwiD83/DSJgibIAkllfo
NFKay2XibdEtlppZtL2z3KIjcrcP6Zrt87YTORqmtlZaO/6oxZWPRfOqHqFm1zFxEiV8w9CIQNMC
8i0IcmP958xDOkE043sjzcKxJv5NILJdVCFecmOYk599nm+QX9MnOObpCnOpsXthooUjNdpGGIzV
OZOpi2HRBspu7d8B/VCQoHMTLvOXZ0m6tANLNElIDXpw4YI33R2n/U3k5pDXwtLuRn/WWxR1kOMn
wcpVSFr4uSNIms8mFSQAFaD9RrsAp6IUedVLwyRmfShH/nBUe27mIt35qMMxsteAv5PApp4QppEH
uoc0w3Viz5qSQ8JkhybfUxJaMRP59HvnUzEeCRcNkw1hzsHrH2TD7LIoBcbV8zdQP+mm205Aep/i
sR9kWSkCbcHsILBi4Yjx/thJuo992oDcMkE4WOn9GrilZQboAE60XF0XL7GIyQmkg+xfvhLe8tUZ
j9m3nm+gy2hg+TsIb7Vs6z/eItgje+liT4H6NlYhpbs0RoerFBq8ISmNGBwxQ2JbLp7WwBeFHa9M
fv7W20CcXa9puu1TM4nWKMeu1TCuJ2vzfrml0uYdbA4XP5bnK18mG6464zrRWIKK/+2Ru8N2Y12/
vHhFpOrCotvwzqe9DNuE7IqctztZIC7Llk0+3m5Pl1Qf073vTHXIYC9F8ZwhQGlZ5qyaCYkNn6Ek
R809QcTXGIxHDHl0C8KqeKKiKDcp0/BQuW8aJQAFVt+aBbVKOGkUDxI2CyjfWWhO0nurJbMRlL6i
9A8aMcrbtoO8gMU1uXkM61ijkbDwct8rHD45FJYCNj9gUa0pPv0PFF6MrywMyRj7qTsyoADO0iJL
Hy/qoZWRhGCUQcRMoF1pTQVsybagGAdctgZrO24O7yv/Kunez3MoaXFp3+IXGqXoWGmPLU4ne3HM
MdyfZGx8+s7U9BE1e6gIm1Mbl2jeXpBErR09JErP4i4AJ5QK8QZSYQzoq/Upziw830sENTnP0sFX
0LtodTMViWTVf2Ful8dwigYbPbycIozUsU/0Jb8LMpchkeBTDz087Pgi0XLJTJ22HgMPYpdR3Evs
MK0B2qHOJQ9mHRNa9V8p8cohBqhm4G+gMgMLwnEsN08v8zvlkv7Zd5QW8HdQlMXzQqvcYbo4q4eb
+OnTFqUguw4hjl2at7CXRn7MDhPxxy53jMSfAR8gk4dEZsDia5genaL41y9SOPfHEO78fLy60+sm
GD92rhO3sGxq/DPihrDYRQkX1waS88yUsqc77SKzVa7T4mq7eytTxPN5d7UElW+uMDs/GVQxmCcQ
upoEEVroNM8N61jtAx5/kzGQ0eK+Gq6ojMp5gm5GB4HEjvcHlDKWzU0mbqUP7kliqIx+jenO34k5
NLOJ35QhqC1LuoabpIR6zRtUYKWYdxj1jxHcgj/rwKDOb8P+zUWuTPRYeKc9vzTMpys0uv9QnrRJ
MOZnt1IdJfCnVx4wy/K1phVVDS1sFQ1nAvfdrULsMxJIvzjqRgcEpWf+yLt5uHZm7yEwIO8aDlSd
xGZZMB/jlbgE5WKfFhKYTc1Mr0a/TgMML3jiyUxXYccXJPWV6tyl4vmfzJJpjB+IzCgJq4i1Sp8j
5y+V3EV+mcjew72H6rRvW0jzTVH7uK9PzMUp2TbrJy0jZWBD2s9da2FCnsDaWYCqdUhkOFb/bRcd
6l+5hoA2flOuM4zSlJIa0p14rh8PMFw78Mms20cIoX70Sjvy9ZcwSvs6O4uHAW42RKMYpgoi930B
zuwtfrwBslZNrSNTHcWNTRXNiYqsN62utPscyu91mZAFoz7DqpoKTqj3g6vOflcCHmWq1uf5enP4
BmNImCL+aPcRQnDEMB9Hf4N1r8ckvOKj/i6v0TR0rG/UQ9AvzF30mso2d0Hz/W5WSf1QpZxSpTQl
sCcF5VpfqTfkpx6ZWRCdLTrf9gKn1m6nKUYskVOELLgB5LS4UMhHRcSPnaEynSlViFUOutBuMwUE
2hrbaG8F2picc0SfzQm2Uav5Sl4eo49K2WYTbQfucS0fWB1pSBn1OVoq7CWPag1wwGJs11+POJwg
Z9xrxLqJyvpMUspHAyZdd/yJhYPrf1sPvas53tOyEiSMAIyx0FAcAnRnrX3b5RfhMLfjuVU+GSM/
3XBeJniuX+171b9IR1ptp19t5qRcdLgcIWvJzmKc/5oHkSy8tofu0J8LFzH5bZO3gjGPiBNG21kJ
Cw/1Jakmm0tYPIlHm+7MJ0kBtDeqNKmG4AR9cg/bKK6xuqblrjzI9Jv1rykCTc08CXMDh+y3KPsh
rdQuj7hA5jX0ZdSmvx7eJUR3/Olqxo7vi1ZbaSKlxJ3G+v68DOeyed1spyGrwfL/QjTr5f0hol8u
eukc4pDfSG6PnBxTuzKdRRQLtxih4IXwgQC/CbHmSmsZZLG9ZWz61TQHDAyxdRPU8aHa18JikDh3
Cyza3nmxDzjfAunV7RAkCxA5E9hZp+oN2gIEz6b8zTdbpqObdTTMlHmzA5ikVodQvNOofsVNj3J2
CbiouE5SSWWZd3S4OznpP3r0LTTWYxA8Gzglbi+kFEE2+A56S1pejkPCl5fuijGMddNBkAKlYotS
0Brt5wBmQx4vpaT886FCkjzCjv6jPzUjix3LxTs0sltiwZihk5U6NZY1T9SoebA6qi9xyqfywnpb
WUCg2PChHhHQV5+82Mhq61dbWLncZiICpR1CejcvbpqYe3E3uFERbTEfgneH4D0ESU9k+gvXu2Ak
rqEDeAkmz1Bz2QZTPZJrfmJOPAAwILTqgne3xi2TXyHuKUNV5ZrX2k0X4qSKT5XLvEF2SvI4VsVp
aE9xZFsXy/cSH8L1qj5c71zJcDZ9hhuaqfx0ycduLwH6fziKe1Vrxia4J/9FHAKeZQ54jV2RYW36
788S7nAYEKFlEW3Fye60MV3fw7jKdeePkuncL91+/f4UzIc7VOtyanYWOf13vz05EwNcl7Z7PXnU
k/sU9AhAGQtbG0nMxnOhm1i5b4L/tCJbx+OaIz6KxkQdde++0sDdEeRE4VZZCOO3S6kK7XXe48Jf
XfLaBFlojeDjhO18rDuG9+f85Ly1Jlo3KObx+ea4M1ulAvErWiTPriOzQZkkMJq/hBLJxLx3G36u
kkxUv+1MasuEjDiMKBXloTKnerN0PXIYkQ+mdDURSHNsh700syLogQEgf1ezzQ6/mnAZQtUfPiID
CcHip/Q12kUys5BnIqHDIYG8Xug/45tbE/Ol+0m0ylQ5Kx0oDXFbqXRf/VGDfwx38PRiBrQTTg/0
YeX85MA4QU2u7jTQkRSAevfCIR8jhFc0MQ7+fbCSYxxtVfyCHEuwM27ILCaQ4Vl+fXzG853PPI5N
V+adxPQSo6sHV3m0nmBzHWuJK+7FBmjUn+wRMDbdAQU496w2dxFeFsZ1qaVbhpELb3lmkvpBC7Rh
tE7Jq8va/VDRoM33ATe1GDs2QvAvphSUREq393bK9/pgvTe82g5wIxbdyWnnSpG9QRWUT56aJPyM
4S+9siqctIJvPeSKhg2JO9t1eDBc2fBu+zDlcGIN0hPzhUOwAQIiI2JLzAV7xMkan+mlr22tf3sK
YlLtm8gvKWrYzE9vLgQJLjIXoXxD1grQFurtmCXdgDocWa15F2DKkwhV6JvSERRJjetAZMbkAAfv
VFQjvbIXGs+c8XipMp0QObdvpgC+okVY8X/hBANov6GESWhVMhHZH2qLfLF2j58cEUXMJL78OA8B
9ob01yxz5JjDdNf9qN+zhSOj/yfpeo/0Z8L5ZfAtwul3p++E2Ys5NZEQyunNjYBidnKHOGA/GUj8
lb3RA0+4MWf/7uX0zsavzNkJ1rfvRQVSSgnbFy7EL53nY0qRE97zIpGlpb/4m9JKx/sdvppCeio0
k1Q/Aal9vePEjQjrABpvUc42qgJP8W+KTbHwrDaB7QQ+sBUkTzMHMSN0pHO8jTk2mKGb88KQ3Vai
lV4WI4kfbEc13fFELSLNsg79kKIEz8Z4zh31g3WbjCk0bwVknTfGSJ91hBGWWbnaT+Jtk4MS0NSg
c5/tF6QC3tEnnMof4KMVuycrj7jxu5ySCFpcSszkcdhptZtPUaNopWA5v1ta6QE6Gh8U2fZ9Ac7U
FjOpkM+dlMDRY3skiaSZanmvvpQztyTnR0CQMILvhMx7Vaq9Bq6GAtgM6vot4NJViN1WiCuN41ew
BMAim63vXSs2Ro4Yv9NMz9fTZSmgMuyJhlxJBa9lnBthYazC0f6xYO6oFmSusiIbD/mfta5Qk4Nv
cGH37h+6JEG4ovEh3qteuW0i6lf0OytWgd3wxpvo0c54hUe7ujWxks+y7CXS6ohfJDcwQnTDjocj
jXtgzUissXpjHxNe6wOabsvFMys/xqg5wW4vcDLW5BZXJFMEdY4lpJHl7A9U7E5Pa8AoNGfnAgwe
vJFlGgKqUkzQwBBcLTwZ/edIxECVOHfcYrnWG1oT8WzDkH4y3LJcHUceSuGreYcjiHH0JoBaAAfN
P80bPhMzGysZ2Z7vgQ0sMnnkoo2P5r8+FvDVVl8WYWZABCyjilqaFei7TX0Pz3T6NKovANoBjh3w
WB1MfDzZm9eW70a2TUWeitMlYv0GRcCyesDOBCfHr9SX25OrXX863YUOUx36rxAuVjQVfDPYu68U
4Hc8hXU98jatnIIPiJvRloLckHsuhLrnx7K5mdU86357pJCB67HylYBeuY5ylF5J5nM42uV0kG9h
x+2RQzCScdWIhcZRD4UKNIryhat30l1T+yC5Abr0G7Brtbx8BGZd/jMNa2T1rKdSj6bXS4rQeUmc
7vvPMZhjlQYE4CL2IXNhppOh9OdWeOfCnVDpl3q1L2XC8AhFbKbq/X4EYnVsHpp2DQrERH9FlrIG
hUUTBs2Ywz/6hQ9yB4q3wy3mRxBFBaKsqskZmqy6kIIsjimFVFlpOq0FnCdcxtpk5kpO88t+Nqc0
C146Z3wioTEVjj9nTcYnQ5jdawJCowrWUd1ygAzPuaEwrGqMHWI1MWlf6yniOkrYsShNa7jjNcwF
t+5zCUi2fbhk1Catfy4vnc7MeGFidJSYZQDE66agWkNUBDMic5wzj149MVWHeVvA3dpdtc7nHQNX
xAi31N9SWvNNyKWZIy+WrPEyuMu+oikENGrsHMsHNXvv1MMxT8SfMjOEnm41ztHP/hLYSXpbIJwp
Y55QOzAspA448fGLqZd2afIWAAQLCh6/penIhMBDqJ+4Ey753D+CXAbeKr3VJ0QPfmG4dUWWZFGr
nCArWGLbyKxiaCMhqeFInunabqpxWdUbMDjmyV0C6cfdWNDa8n2ARAx0xiG3zuCsyFrsUoxsWsbl
9mlT75r5RJHcHds+nGTdmcEPf0SMsq0YshedRrq3H9+3VNVjOOmi1kcR22gjqbF3uyDWjjnO3mFp
IJU4AiaUkOlTIus5ZXEKoDohM+1WEWSg+laFFyTR2YNhs/96OZNxBmYQsKV0U4hjH05n7nwPP5Wa
34kORV6SoJysBFevkAEfHeG6TIy8G08AcrXbqswU06V62OG/BxIaL6X46maZ6nVGKqjot2JQCwAq
r2KwyNXZzSCDmuD2AHAl6cuXPDbBWR8V+UkTyDJ/5LzjS8nviwXmh3nM+IDAHqa3zXHXImPXv5/K
OG9Bk5TJR8F4Y0iXAkyNV5kGsX2MRFoamsrFGOb/QRqNnnpGb6FEglmWNphldNWUqwOaBMp3w4t1
j771eO7c3LNCbhO2q4zEN18KVxb7al04nO8g6nFpYcYphFOifnMlqno9Ui5ictX6pXgGXrQXFhYr
I5UKZfXm7GATqjjzAjAX7WZ1YNKCUuVSZwrMUsHNghwqOXDQJ7VKyTGfaxivdTTW3Fqwu5356UUH
ZLg5wHZO7h168nc+JFLsfTo3DXYVweted/P6i520+69ArE2trv+YJdHKT+2NVA6wlF2/i1uFVQBb
Jvsk9Jtt/xWGWDt+OJVR5kOG9xap5V0EgrKdn2DHPyaFrlFlmMwQiEC3++vdgDQBJYU0YUEKYUyg
cKpgj9XXVJ/mT51mzdmcqpGCTBcWfvB/s9DzVFJlE558jUzgpipmffKA2T333suxPyMekz+7i0B7
ZXvAcREoY4btTRkCTpw6NqG9iHpEXUpI6w7pQiPDXOrG8hlD0fBNutiFcxSGQzlxhoQV+NTqXtTf
Dfmle3U0GSV0Ocgdhut6HFgFq4X9448UxM0Fn0spbiqSQ6glSot5P2gu07Kq5zshxXmXMe5XCF1S
SWSQW7AbEickwDoZ6Re2UHDPXEYiW5TGgiQnlYbH/oECZdPL/WYJ6kZF3wNnRvvUmN8kbvrXd9np
H8oblNTD5rBxPfAueR8LA7QcAmQ2oiQB8ETWQQeLvIid8p9ibIOgo19sGef6hQSkfKPESguiZrQ5
n8/1eqF04aYNFghOxy5DrlXgrlHTJraKaufzEdOu++qjksY4vkd94dGMaSisZd36hQuq2KI7K+UK
98sE/AWAROkuR4XlWq4KvskTWLNhqwHGdjvAb//XSN6T3yNXT3udJufjGrKrjN8N7zPNKUTS1t22
jvLfF3br5y5fB4k9hhtUJO7UYfoZMYkto231bKZoUyageK/MqzMSIsEwCoG4R1z8lgXy2ZNm+Xqw
MWZzOf3A443Dp21meLULGFLhakAW36GtWz72Uyu7B1zGN0c5N9fsyyKCieBHf12wdHSW0qUL4s0+
8/kknVFTFMLlp3K0b2pvryP1Q9s8Gmf84rOPdB55/Hm4iYzJW1tjMAJ2aXgWBXcQLtfmhoM0eIB/
YMwgiIGC4z5WUsmMQiiIhDHTrFlHTs5QvDyePt3e15Mh+EG8KN+XoS6qQD7yZlHCdJrQyT3tuPiC
7VrVmfkj/X9awfWlEuIJ8b6qFr3SQeaiL7plCY8E2HRkp45MSKKoX1cvpzpqvy799LEdSHpx8IvM
l9swRy9YC3LJ8SevbkT+IKQGrEmMTlo3QuERHhOdi5MNqEtrdOnQE7fCWhv6uYUA3qSU8ifuAT34
jbtRO1atiS01gx473uK55X5J/6ZykCmHUDxNSI6Oon8IddsagsJ8PVsZ0gsRlF0P/HvG4LB5bqkJ
KkFkRThtopLtJ4N5H1hiTnWZeB1kFHNZZ9mLx1WnYoxSFYSzmqELVy/+zdidqA5oHLpWtwQ2zBWw
18hFoPfTAWcwCE6rO+ZcVAZxWosyG2ZWPLxShQM/zOU75WTaEw69XzG6ZE/IBKwDr1yPGlbuJgKj
MSF7q5wOtZZYQ5rOnfmFrWVs3Zk4Ky9+bVtKf3xIxttxmcQjWtTrB5qHY+bQSE7oAUGsaklMOC5E
ksWeaB+icnz8XfAUbZ+a9PYq18HaRb9tS6/2ZrHVOnshD54HSPgYfQ8dS4wuzwPqum/V5R1A3nG+
vwx1/VUE/YzWljAyLtf9Xl5pFtg0nJ2kkFj0BBx0aIGOAwQLJ0OC8LBTxGt3/FdhT0uiop0g7gAv
j3pDdP/ZFUJabg5mDHDa6eNxF9RjLw+ncjNr2QKGlWPna30qm4xa6jyCLom+PdotE2sCKWI8m8X7
ffBxjpAoZt9JGKjolL0JIzGLaf+d+2AsRD8N+sHcl6kwvTcJbjx80w6wwCnivzAf8RzJaSQ2rvLp
1gjNZMAQ9+KUGNs9ThFiaw5nypmAE+dkyUiRmk8MdbuOeCCmRxbRSUsNeFw9DyeI6OzBCj8H2/h1
imcet594uf/538iEsvygw/UugdeMv7Q9bvWSEVZ0Y/GIVtLSdrdRYfH2DeL0wPhME/LNgUhst0jx
oa0usuA8obWImCrCrS8JGYVMMAkitzGtfiouiOBD21c1KLxJDMyzCIxviToZYAVcj8vZoAVZER4C
kqhWpylVi19WXeLwarvB92PRG3utMF6Z/Pp70p/yM6yZBSVIr34WLiJz2G1NQN+DTwrk702RF5sB
qjBBUyO7mP/HRb6cGWZ6q2lCtm1cZYkEC1MkPJoCwzP2gquByBvzQynMOeFkXdqizO8QBFHpBEAk
rinkGtUUXP7cVNQIwXgSbBN9e1u+tgbI74In4XrqqvUFbizdTtr9qY+Iaa9A/0gh6dPkYN2yavbz
zIrUSZMpfhpDTm2G5NQXdDP5dtR5YooLzcgk0OyLXb/eoFlprXtoE+wTCq9NiDitNVWi9gw6e0KC
72ZMVKuRULtg2oVDXkiHuoJtp1ITDrRrq8l8sdOwlcpeBX711sY+dvKy+IxqhrCRQjY6UhQBzuKA
j38z05lYWFWmApBOYqeXHWu3cxS/L2OcNk1+4YQLGRTMCs37hcocMUC0FO1bxw5ysVLHIx3yuBRP
9wJApgZYHWF6o2IAzxxxXJpqfe3ZMqEY8d5Q1oIjXnIMIbSLD2a6FSI/McDau2HmiDEa2Tj9BwKx
4VINJsTT+Q6JZL9zqxYXmSgNEfRtd/HUFgre+ojgELH2bnuF9Bap1zs8YCVjiN1hUrHF72f5QUrF
jGHxSANK6nvrqs06J3qg2ZszXZB0QZ96eaUtB0+eI1ZMS4S+N1UM27SEbrCISi4zIoMTnJ1RSQnP
vjU3M7LduY+5Y2gQFCTCvj/ugGK7UdKaC36TuaYnTKsnHO7wkiGLWWNtTdy2lRJk+0zb3GqzEXUg
a1cPrxnodSuT2yRzVq8PqqKortjCFAWBnjBsZw498mp+55wt6U+qJ6z3lh/FNATL659Hvd0mKzLY
X1iF3g1YAVrETcHnPqS7q49gwN7csy0EfBpTX/RgHvZSdIdKvc9XmxiUYk/dBMXh12w7WH8Oye3x
VEMl6bn3ESBBLaatPR7MBl22VDwuQ20CM9Nhkjx+cqNIOnUgiJeDUKXmDesHyOjpzptQ0WKO3v09
udv+60dqn+rOPGePrITNaFbZoOWDwtiWctpmhaZbTpizQqsrzPm0tlBmB2Xj66RV7W6xhEzUmyue
O7/+ZC2B9p05E7wHs577RDx///8Y+LHmRgnQDLWE0RNPmama/q4Z6wxm6OFhUjXgJoMt7EjYMrbo
tpwQfXwSXdZ7eAa3EAJjz8S8yebtvRFI60HSnETJzPKxtjussX7Cp8ZCMwq75p/dPQLDQ9WCQEqD
cno9kqx7pNH6uhYxZfWCuYIgn2jNCkVLnFaGoH9uI09vP+Zwn0QvaVtv7hJ+MLMpljb5yGKxARVk
K1n/aZhzd2mDGyXQfKQgxmpty/Q5jvW9ufXaQxZ0YJlaJyOFgPOaxuL5uBgQc6Iero37YArWG4xF
vajw1dkgNLDxPkbkliog2THcozh21lM20/LXZBLMV3KRBu5dktH832v/5XDU/3MFWSZEunUqpiOV
WYYAjOfhDSUF1MeqP80harhUid+JDfV8PC/4wg0ySr8nfAkoRAHkwfwFAfgZCB3tIUP6oWyljnDm
A8/O39kiFrUu9Mv/cqsh/Dg0LmeAzNjez+NdzvR5/wkSl1Kj/boXCncZfNEYyzaeOmE+fTdTCCMO
FV6Q97C4Z5pCWMyVMDEwpCiht5K4CwGemW1/+U/kA3y9G8BVqqhtfvAufgwVnSsNkNnku2bShSds
RJZqCWZCt0blPj3FLwAOmg6KdItkLwJUNluuzur+JyMDhBPrL4oF2lRDpOH6cUITbavGgTdCougD
OvYu4ixZPJeehRKZMur+cC0kMx8aXPRMxxztjEX7NTcJ+jG9tIyZbpPbKrVKqVzr+SrMJjTfgpRH
lv6BS+Yw/hb0ECk0v2c0lzrks4pB/L9KJ+XGBADAO4ki/JEkDlJBq8qk99KSXhxvUQqMziwaPTZh
KZaS/Ig/78VdgPvULvrPA7p2FggRa0z9HpS9H05zQPJpx7xM7LFaDgO0iVVLMw/Bf2pnn7XRO6xP
KQ0WxphOE8Rk2VaNJQYjA1LxkyeSVaXlUX7wBCJtHwQBR0VZ9mxTfMMRwxhvPm9pHLThmKMUXQgY
ya9Pnr8QmnOUnIioPiK0EZxgDHS+UypfJEdXxlrjfMxW8WfoZC9qGdNBIGZiiIVRTou7FjutUEBJ
0gFreL0DLv7I1ZBR6Nh/V189Z26PlIGd1FK8jf/mYUe1O10j+yYjUT9pEtgTu1E8ZXJ7guuUL1So
XvDUc5qavXg07vzGa05tljzADm7CxSDWkkBhV59Aj1lBaKhW78+pMrvw/o5ZRAerA129xtYBKWOD
FgHt1FGQNTPx/jU9C9P9WWdeIcWcsbcAs/wePBkHz0fX5tHtzlI1ltU7Z2BB0+S0b67/s64lxljz
X/WTF/zeizE9eM1MM2ERRgoR0JnzA5h8Ry2oSL2CQDf1CPQIe+OpXk6BQi9h2u7R0aPNFuJjcTIe
QzvuI1pPO9s3L5P3gO1MytS2i9vS3GyQjjHCDQ9cqCVJhNeJiBTVj7uSGyomguER00Uf9mFnw0ni
1znTzu0p2VvXh44I+itZU09uZ3GbYDYMznONWGnANDnfZDicdA8YNx5MeHnzL0YqlMCLu000XKSw
nJVac55oOQYJ9qnMCqvHvGdzZrAycNne+yfUi0X76TxycQdWR0h5AQSX9Uf3QJ2016cjhF2nRQhV
YeY2sWkbe+0AB6F5U/wGkI3TaZtkbqiKXCZg4RSOTxXvy+ctgn8a7tzGcWNmLDgGqePdml0Q99Sl
BgF9lX5PN4Wms8WbvJeVM+iG/P6Wcqakzgc5f0SIMgSfOFrRvPvwo8tG8udLGBa6jpyVw4sMRDVo
D2wND83aK6tsFiXo4MV7hq/WMy0eKDKQpzlTU0RYMFT5OaMPT5bMBhOyniHYZU2gP8qrxS35bw9B
EHq+j6foAxFl0tCOMnafjpDVbZnRn7hjBYFQ44MH2a9uEeSttXdfwwIBzaiRi4g7VsKBC1HmbKUi
wnDUcb1yJhmPEBSEWx5mCRUvmhhBbg2T2hulp6Fhe8Jbi8I0wt5ohhcrxHurXuXYCeYMTxP4HmaY
W8sPrrHjGKGS/GevIP6idK4aebR6+uP5HzvqZynQ/1XVH/J3H1k+kGEXfiR3MDVnpRRpgL2GRz13
0llLp5o7uELvtw+Rn2m9RN36qlkfOfb4cq6t/8SBXIPR2TKjfEny0v9I7Q23aoNMVWD1xgO1ObNH
GcYgN9UqfzH/03+pZ/CloJK1Bk/zDhxGONWGY3QuYVU3TfSIDBMGguc4VKX5MLzASsN9JllP+9YX
fq/sdSt537mvRNXHnGWxkEaE4kriB+AIdv/8mMpLTdR2UmQB1quG+LGIVVWZQjL1S6GsnvjfYxd5
ug/ys2376KqpvCowOSCXnwoHTLfmt9gLsxIg8VocAgKVP9EmkilGS34p0S2sc+sRSPYYrpIXRHRf
FJZXy0m9JDc6hJACRX3H9YmJ1X/1aCG70b/06fdipQ6mhazpv14FiS0sznlMA0piBBs254GBhe12
mElDdezbP+R51cTz3wVz8OyTKpA3SrH9nGA1DbqMZGU0MEE2B6E8+vgHe3MCMCRn69m56CCAIrNR
2qU8+jSYUdfmT2a8AyMiWUR3rNaR5LPIr9ky7sDdneU35oBgO9WG8FOsRLyWqxiS5ZLoJlqVIiwy
vMMqPT+YD2D4uE2UFNf5NsIPwosmYUzGxzU7QHKFq9HCekvdJbb5VPLNP3UJiBluBsc7ixl9+RnB
VxIcfO32DV56QTLcd42XPFJMCuHROs0IHiYNXbq3zfsix4Zn5pBD/wRDGi65GYVhs4/Nk25WOJ9g
ElUerbfLMNjxmI7i7TI6755AJlLuhDptMJ3pxB5EhaVi3Wr42fw+IPWWbOxQlDwW4sD5D5I3LAAN
FZ7PoTzZA5u8JIwFtIr7ECjgoMzWLXoSfyal4Vb5u4Y7xzMt/v78Qwwfjdwblfekx2wNpUV3mJx6
4SLx0Q3BN+hsDXNtK9Bv6arKQ6qCE9k1OVR+9HiM07UNC4+5VYRMCv0qk9kGL/bZGLVB2VStVuwp
MxaNNH1aKkNkYiW2T4+ocM5rSJSqjFOWv8qJyDSb3cEZJo4QRF47RqRcGU3HbNXiEvvapANqJLNw
GCPR/PxdMYTTc3QDZgTW49SQ7gc0pZ4bK6elwAUAOaIVDSuDjop7yNz6xeIK63ymjUAtDkqiCJPO
nRGeSM/pWXFN6QZka3olPvs0lyi9JeHeYD/t3Y1e9Jgzi1DX6n+o34rp8po8pTQHKWPPtPMTcOHm
xnPs2bEmnsvl777rJZ0Bhls86tdmILXefusgCjAy8mb0uQNDpdak2EkwkgtyakyBl1a0YXvnmzD/
2ekgT7JvkBn1ze8w9CTi6fkN89GnNQb8C5GZiAO7KLGFMk2EJwkx0pKBu22ch7ArRXYVHtoergK9
lifwjd0xTBgfv9kwZw6/X1MbZ+AC2KMVgCQxDCDs5B606W/rP2ETz4kAsjjqL2/zxXKLSCgUZQfA
jci+cOB0BkzN4ANwstVY6+Qn6n2OprSWsUVjOSzME6wJ4ZDyswvcgbld++NeXFEGABWBmP1EwPc2
E1SfmpmsYXA3iArR4q2S4uskZmL5mE2BYR+Sd3J2g6YFeg4nfxtm8ie5Q10VOKWIuCRutaGFKikb
o+aFfFA2vr9pK/EyGQn22JY2FiOJet3sDidHxTSsM9Xr6eE/QZpDsAhAI93q3uLyThOPlkmW5G8n
09L9HXQGMMDhgSnwuq2maZTNZ8t4ixzcvWdsu+BJ2kDUKIdu61Tr3fnd3n/UZ0a6Lzo7K7481gCE
1BAyHVisWMjz/7iDVC+Nrp8eilQzNC+f2/+Joc4pzpALBjmDwPsGJR7UjlEzJ67Og4NXXanClyX9
aqB6ZHEpQsBEbkNaWhNAQ6XGOJN4VnM8sgjJljMA8+nwVZR6nfS+PHPT8/Cq+a1j8jjQSZSqw+C6
MWIjY2j2gQ4zejezjMuJgLwMoE67OvJogyDLlWyQW14OxLFW1qjne+vEosq4lOeOEP9EUB/2/kON
02LgutMTPhwGEDG7XQY/fQJrhbIU9kwtHNo25vNAPb93jzDX3AHhSBAxL9wmWg+CZEoZyOakv0Fv
hDNd8txb+hh3G2bfTjSou6G70mcnYEDydXX4NJSPn7QhiL9JxvGsy9ciSoUe4zPD+tL44pT3Pizs
+1D8wwkdMZiJ670qNdLTbYwQxoS61EfRUv1EEgviQkKzJc0WbEluTQlaoUS6AHDot7L/yDnZEFoe
bhAJE85du0rq7BSlQ0l4WV63nv96gzR6hlTcQjrE0c0Jll9VDYsiYeFmRHf6DLQvhb7se8hYw3T1
MfqWr5FlqUJGnLzcVLDHjy54Oc0WENZo2wuMkGo0F73EErD/aEy19wLj/auOVWVDHFPtXDBaNYZF
6l4U1BhnBiZisDroogSwvXoZTswMi+sCdsq8VFstpDRb7eoXLLc9zuUydbv1ItvYgnbqVtQVC8nq
55+i7cB8wEE31Sdxi6yyDg34v0N4nYXGe7ymWfxs6tzdxQg3HzIaOLYiEvBNv+9XqtWtyoxqk+QY
rqJHlWXaZVMWNPOZap9Y66tjBAHS54nFG0fUpej49Yc20OBfKOvvaYmqSw0hbwrI5XJp+WKr9Sp9
f0B1Y2AkBNxTBZhpaoc7RXLsWmWJOWojjaqM8n0MDVylxD+A3mdKvmBXP/QhHnEp8GRk1ZjW1C9T
nJlabBH3F/cGhPulpJCNrXJ+oMh27uA36HBo3+EpYh09/s3VyFKnjR8vHXikupXGXsDuCDnil3i8
jy8JwMwYxC7CiMW+aQ211covg6pVEkVqIENtNNslUSUnYeZUesCQpYVBWebmLd1/wIr6oj3E4bc/
5a/Qy87/egTge5leeK1G6SIijKVJrXKEYm6be4Sn9LwleIpexsENAigqsjG3eZTnikUtlPStYDaU
hJS/uGX37fQk2ejUxp9Xngms9cDSosfKVdLXsqqrjjqW+3fO+jtRHT+qJwyhFk1zdl5yCQrHW9VQ
B1O/b1UgAjUDgeoRp8QMBAPXmnXdw/H+CaV7IjrVsAuO05H/kpEF3oHJsk2fEecfxSNE7x3nUpt3
iJyls16O6I6edfqv518KTJTpMKwu+CnTCXGAecNMvN8a0JI7NflDeCUVm0SNujNY2uz+xRzbazXo
3YZit8SwK71NNpxoZNCEYaq1/g5JS6YqQF/EI+ZKfOjVp16d0Gsi/c4lb6BXsvJi9QYCugLIgV3n
EMKRMou5IvDQVUp3Y6uk/tsuXXa6r9eA9u4ReNc6lntMYuXbIuv9QxF+cmvn0SPG/KfL93qCO50t
LHj9d3YGudh2vTfx0r03Cm78bU2CgU8H5b/tDKKZXtUuPoa++nerBrQepgmcgJzdnRx+dep7MCbl
sIpTMruHQXkYO0qHrhPKxT8gfZUqZb0zj3jqxeVSZZNujGIsWGcTz86P6XJcCmZmQc4G0XtqtxY3
eBe9KGJIJEpukeaMZizSzMfTkPV8pNJyF5dWZRRjKtc/idGja5bhXAJjL9hYry7kXCj8ZrxXyTYd
BvdbSkfURXH0RJsjbunmvN/9BM/UZFWBM+lJm59d62+GQEbkxBfRxOxELwaT/YtHjc9TIZckrKVs
rNAaYC234ScjVsD3k8Hk4ywYWE8aiTPV+Bh3Azp8nptiCWjoxEWwlzk2Zbc6qg/98JM3rzExDBGr
jojApbIgW+H7JLtCmvZILqT4Wp79ih61wPpRtBVnbNTVwDLrRphN/0NpEEWqMFqmJ7/Jvtqb2WSF
spYQN56HGuVBneXMzzSvAbCjU9Kc+iSYq1VIGpMvwICIr/DHXkWXFpfqv8+COmAul7ljMtog4m5h
wUUqloJYUHQvGF6EHZN6vpr1hYxFvYYzyRSZ2bFRktWWRykqq/BAOOJD8cl+36tt/FN8Wv4OZnI2
C9L2M1oBjngn5iWTYaBEvTVAHUHPB1tCeHUd/ABVqTFJnSYa6mIkXxlG0ejOkFaUEGs8laPhduLj
lvZG+mzFOm5ac016y1Q2R070b9RWcR/AiwQQ52+gdzSL1XPhOeNCWh6+Vx1pq1HHO6AufwZ9WCAZ
VZ0CZu/3aTn5m+RsNuuZ8/t69kVLqerqEcVv9kbXp5ImufhzMp/k1YhfvIecAcATy7lusBbVbe2G
dQpf2IQ5YIEFKcF8DnlesaHa6DmCYXGgvrnh0cwUZhATpSqT64iEGTkSrsmm9wBzNNJHNXCzFZ9Q
FbeQkdszH8dSf1AuR61j5+zSw9gPf4U0ZLxORrP12vuFObUg7hKKEpweXJ1u9xpikkJIqHYhn4GN
apxloN9e/rnf1hRF8oh60nwCzillu1lUWhRsejtNaUwexgDTszNqGqXzZ53cHRtdv9dpXRC6svsK
39i5C+pSw8zTzBQPBe8a7PMfHYMfbUpiXWVA0JcaCaciC1r7QwwKXqGmX1tLddtt1kkrHYGvzP4c
NMSOexbqpQVQyO8+QLMUmC3hKdd3lb8B7A5/C7l9EiC44gQyMAR5v3pz2BzSP+SwYiRexckVKaEb
A/0xdUq2wLD4Ho68qbNamrZ6tAaQEhjwnXUjJU/KOkS5hphIGHBtHRDg/cSdtzJ3ZEBgx4nJIYCs
q8F9DlyGh3Tq5QAKeW+FxrakrOmtKNymL7ihlihdXmD0DdoxQd0ZAmwLlUpiSIng320z6WUE6HJp
pL4JKV7PMxvVCEV/R39ZdqJhxBT5biQqvdN+k5rmZNp1FYvIT6VBYZ3uGV1fjK5aos7MkEAAdR6N
00n8l9RDsK1n+sGHpUzXioj8iCE0w/xuTIJysfwqmR7QSF85YEG41mIe5+YfSY94qfE+KS+oc4LW
lhAaa5xYMXdjcXK+1Ng1WWQQealmMR7JhkEvuRc+shVadEMvtrgRsYWrGgUYbGduI0YaKc61B0S2
4hu6DEy1RU6h43/rqZc/RiYi3SmmRQo9nEjQ1SC4GMCldotKJi++1cpgHmhz8tXIa93lIv2r51rV
6l5deSTh6989/St893C4vejtTKDR8r89//x/utXdOqaif2EpQWsMuPhBZpVzSRHUMaKJTRmb1rOh
rU9OcnBlAMJggFubJlAZMnxDA21HB4S3xgS3+LEqLYAMmOWIkyLavMR8QXgn5FBD7F3mnd75w1Dg
0NH2v5wUXtq0ZMhBlNtW2cAQdNzkp7siexuiNjWH8dP9avxanMwdrDLreO0+oaiV99ZH7fGBn5/c
crLdqi3ZqDV7wie2rmp0cP310/HIJOoxeQbcy46RAAr+/64a8AHiODLk+ikk7x4Af35vsXHpnihb
BvtpeCJuEQByw4bX1KgnFKUqg7FimzLIu3nufAUybkdqiYZSG66ziLqq9vgy8ULGxafwxLoW4q27
BKpCDgE3H68YBgUwp0F12Ho4pp7kYvFbcltY4fNSrEczXilLeaZJEKEJ0UCgowfae6mDCvkYwyrz
Zk6lWqNpBzD9irqJb6OBnmH1LhkldDEGxxmjPUJDr9CFK2eQflqNSWchdpfQCO/yuVW4lMUolMYY
Z1I4Hy/HSyddF72Oep6nLSK6AF//UXfIf0bARt0Qjc0Kepb13ClroETCl+J/kF1b+sEeEFoiZJ+O
Zk24KE1iUSN9iclfOehSccVyrbbuG2OC5KGCV993eKkmV+cMg5NxmPpZWtQh3FKdnvZITaOSi6Ov
UmEIUUYYgszZqhmJB4aJw+Qwg4daQTiaQL7+LqylZA2O/vnM+fceC/JtnaHMvKfJnD6Vzc+5Rd4y
EOLf/euJ9V953/F8weJ9yNau7C4/Bv/opTzQqe+s5lD3v+QwX5iSubm1zMIXXztAI7ZMJVhZ7l2U
AgWDwM7iYTdU5YSEXdVwUJ4kwfHJt+GauuKDI2zW8vARv8dEeUvlSAlbhFFLAtJuNXt5EXhTubxb
NYakJ4I4DKFcxnfn3+s7Sf+AA7tqDpKn2BJgjdL0X0Y1ZVTYov5qnLpZ2nSu/ovWucYsasncouI0
20TMeTHwUAdhGZKweDbc3HN51ZQEwX/VvV+br60e8UagMsJJV360mDwohnBEsRMMNxsQXON+LXOH
EsACukRnWpX/lrftNJaH++w9wldcosg3iDT//+NErBQn0A0sR90O0N9toTfnjpembWmQ6RyZCjH6
yNMyFWvKGAiT0Wh8y4bhkejK5PNJhK3tjMHE9brZUp6YZSzaS4d1/0ZzVUXtKakgSj4CYmIaZHXQ
QFOLC3gWpTnw4J1SIUty3oSqaCH77BBbFDo/WBQutdYkoVzVYjN9kvzg7lzR+NuL2ZAaCyHr1uiX
HSDXm7Vnzg0EYFt/SxrdaVtNiQVzSjcN1bsphlTc0ywEzWebOeasE+nyFYiLoWqNUX6wfSr+bnpV
ZG2sDvHev3nhJ1ZOdyRf7tDI/qq462x8NyePo5yrzTvSnehO48SNkAuqDiZgQLeNr+h8aj7diE5o
/HGMTlz6mcK/6T1KiQ+QXDJEvDHn8CnFvC2FHT5/xsUzJV+DWcmrwE80sta4SDT6Irr06GcZQVTk
glVdjhSKe8d9CvmjOuIABwzjC/B6QYy13345j+uHdfH/xvtRDQh4rzyXEcVexNKUK5l4JN7LRvPk
JhUyrJeTaWw9rUAHoZD36NwQmsZHXQ0SBDeP40QaBOHvSF6Ea7aevrLh/ZvzSyY/iTfr0r0q+tjw
HCtvTsURGlosjRmfitDlVfl5bl/dUMYfhVk1JAYyNaaKpMYbgvA2ft/Q+1srISOeWdeFcimGF1yC
AECeZ3L4afN/NHXBlK/PdturIbrTMyAbCuUAifr4/KMPX8HusjB1TIjwX7ulj9UeYvTYBytUtSby
sGvIC5Ri0j7LnmbzOYsMPRxrOXKefuYfZ/ZHpMjAz95MLrZk+mS+4JYk2zsOp+Jdmglz69kMm/qq
uD+Nmqm/1bDdbt9M5+s1iGsUUHde3RytmAhuNBc+rZtdCoDgEZER4HOA1HM05rQ0ZRgiSun5R3oz
vaCPKujwZ6RbclVoEv65ZAUIH4heq2ElPmIJ+77VVZ7PP5K/XZNOhEFOSj6302ydR0AmIxWbqAhN
8Llg/JnZhIeMUbPBhq8ATXtfRVqU8I7L91GTmZlptvius/YjKR7mbn2k65fMy9XdVkS2NH+fGBh6
gZm8+od2WhuWADK/EXyxuvNpnJ3wbNh4/qsofCnpd2E2FVSbncPu1AEyx+7z/P0P0eRwiTmHFj8m
LfL2reFF4J7OjP9YXQlu4nV/f/ftD3vw0CnghgVCWQFJWhu79RTG6pQamzsiNF0cGbsYJBboMktP
z7K5fLhl/X3J9iuiEwtHRF0HQWUbvcv/XI74NtUj+2pYm2ehnv3e0GTJK+eDNenJVGAUaAmwNnnX
eALpBbipfk3iQZSGpxfaOeYhBPjmDbwPZ4vlRd+mAcIZlu4exjSnKpM4RBGRvV7xDCNy30/AvD+b
8VKytVChdSjBo8ETvsqhzwz7IOFuPoD97cvROWtBbqC7/gcv4XIA94xgI/Aedm4MT5AICdwja1p5
UQF1M0PfwzIM4uttehjoM2YfF9Ci6PG3vT09ueEJtlzXhEZgyYuSnCeoohbz+zpzfR+7xvviZW2A
rHZhUcHgU5bpsesAKpZjvggZl0yTNNq9C+4EYCVmKi6P0Wgc5mq+jB6JK54N+8XZ7Wn34faUdlUF
RuhfRnJ5s3CK0qWUGkF14oTxZSEmBjoH82vm/CR6iggMjBiEpvPX0qh6j81g3LV3FassoFds55Z7
rmWDCSZtiD91PDydqZRnDyVmvleVgDTtBeR6Tm+x0h2wpOQbRc+juz8dJyFDXAEhv9vW+8oD8qHa
mtW22WY/x75RRjmOI19LuN2fYleEwxMyWPrpJozvn75pVSeuagpDZaGL9Y6xzO2BpnI8OaBt+Jae
94+fIQFAwHmy1Q38sectsRtiB0+SVQwp0/kPiN9dR7FDIi80INlzuJqvtnMgKsyJ+QyJFlvGDnI6
42wayRxL8871EmDQDCZY/nka+9NQUjrhgey6M4XXngzkbioqLLmF+Nwc8QwuHp9aZNtoLBooU6Ja
eWoHFdCA9fKW16H6ODYXNJUYdCdLshw2RLi6gfoqZ3ctCK0TGqht/YUem4g+XWXbwISiDbVqjluL
cevskXardX9QXZ9hHsfHbNT1FviDECXtlhXkUEGFPbjMRKeJzaIWd7sh11jzphBzXs6z1D6NNU5S
ia65rZQRYTBM01krcwqQCQR9cITyD5VgxIGbdwsHxaH/GOWedHAnOoolAIfj/Vi0SILx4bd8aNwR
qa+mDo/2FxvPDGVPlxvEVz5M3jYLLKuSpVrDa/sstXWwSX3ja1ZLKGUEqzHqm+N96MJ6D9NdH5yl
iiVWyDRlGhSKvXjGamvOMjv1o2QK1g5iod5AJ3zGVjvi5aJSU38Lbq/C6UK7HEV4cAI2k2jrScy6
oPdhOYeJ0MsyDtktvz5uqRGqWfVIhx3Lhts1krByu4N1CyVzzYJqc/gXVmoP1wjDJFAcYsg20DWj
NA+OY6Yp/HXjzILh26licme01XoynzblEZNJPCL9BLJoyYu5Cbe1ObW/47WHrfDlEq3ciSXRtIUl
XCb0q/I1KXKZvjF6AYw36EEK3nnmoI18JZWUhTvuRvB87olQ2SrOBlW7RUdYUh+wc8BgCKPj7PFr
LVxzl5Sgv4b5SjzjKUqVySC0EOkQmhvH+LtunEBzLmkmbSZ3tNGAWEAokTQg1utk0SsA8OIWBNWV
kX8anivm65P+aIe/PRB8zG1PaFrZPMtCXPh1lE6QrFlrBNHgGjl26t57zga3T70DWKxMDcL+G1sv
4zWOOuaM3DhZ6K+9wMu/9j9RRu5lzzDW6tLR99uAmnfJ4bElQzQHvvqzJ7a96wjRfkp0LVva/8Bf
1bklLe6y0nhR/OYBl4hX+bzh9sRGLnI+CurDudkCSU9NqZsGODkmqwu8HP+RU0qqbeWugy11HzZT
G2bqxQPII7EtMI+OgLXfsG2x3P6ihw6RpSReZCxK3U3YQ5vFq+qgfN3X52P8z5ewUfv+U8HEJHUp
CpPY91oSNytlnHrCJXF+WMNnafaEnxZ8sHgPt+aXeh5lgK7DX1FP9dAT4Zg0ppirMozpp/kqYZJ1
VeZapDyLYtKQfB00igG6a4TIr1miPCVa4pW7R1ymNAeLZxcMtnMxoWlZfmnp2RyvJFrmD5aS8kW2
smclRaUrYzg3Th9LvXk1wKCCAryVQs86B00KhopBYgdIv2k/BRxlzpN5RFlaxw+cNMdhtURvkljb
os+lzpKj69lZt2Hng8iZLVIW6kLIQfgW9J3A9PAs8j5bY72lGFs/c40hKPVttPSMO/3arweto+1o
PnuG2GL9UO96sv4tNXxEkxXN2DVnuOpDv/FIGvG/jaV7V1586v/3pLapwn1IC8yeAMRqrsnJURS3
LXsij3mQvCfNcQbuBlCQl3AqJ5nXICDtWWj8dUbt9TaoI/PilQw7sKg1Osd+LPN0m8hVzvak+VTi
0k351EbmVXFRxI6yB2csZraBHnVixCUiA5Xkb9g2TSxN9sm/RkVsrEG1OyqcOC+OyemTUp593pOb
Bx36QbhCDTjalfM/HSEnr1ncGtcwlB1XtkizsfW4eJ6k+kFZNSVCdJALAhFvuXw9a0E5Lb2NrUmu
J57JwgUdyimRkYLcRg5cqJZF9S9OYvEhvZ6Xdms4M7/9qHFeGZY7Fo0EQg4OWlHkC5iFrUejDs0k
Cc8/PJkIJLZJuqz3QoO4c/pww6hjTyuvHCiNeGWCjK6qadV7l1HImcu8R10eqmHrW4Ar2ZALV0BN
Sp9KXiGbS1Jh2kiZ4Y+2LZ3XAVBcJTbSRwUbfXxJl+3qm3g5Z4dipR/x7799up049eqVzvJOrjP3
ewV3eWCNiOldgRuRVtd+rkoy2GC9V1J0VooaKHHmfV+gU7Llc3cdxUKAjh6WBZkpCT452rt9Hcws
Un7fxQhLubGUm2mQn+quboERhlaUf2GgSfqp9ZD9TDEpg50gFHI9luaUq8GlEHpYER+xdGU4VF89
HMi9UxCZGhVnz5/YzR9g9bpUE//OwSUOrKTN4y6XD3NeFzneVWmUrKDecgP1DmdbpbvhtZenuwgJ
UsG90AmYMZy4WZQnBqgbxLrkOHoOz5wiYfYkxo4uP7KUhircYYeHQMS0+34BSCA+R6uLGhmdIhwk
jOq//q1peWQsk6xT+lOpR0dKqCMOpTF4fk8C5pKRI2ij8/5mbRSQr0zi81KPaQgcFlAv+AkPS3ZJ
azVwlnqwAUxNxRSRYj+D1f4eYRMt4RKux3KJKP3KLfB0h/X3c6QdAyfNnwhEXUWDFY/q3em6Kbm+
fzqlwVdU+nr0lbXaEmsAVve3acH0K56cjScaHGQfrK+zr/eTl8p9kLEXXCl0eUEKp9rHiFRpdH2V
cOgUfxrjqfseLIjQvC81NNzC173i/zEbjGa9pTITgD0cQJ1Vz5fJY4SAZRlM13CQdqqDQpHzgw08
qAuXzn+JgwvMvlF7JpObq+H5t2ZD2TFhtSYFXekWcbFZbX3OuFPWXDwTZbz5IVDMJnM/i5WzRhI7
mWsVlOr3sKJaHd4XPYPWmXBCdb+OuHyXR95jzZQjvA6FsyZh1FjPZdGG9KfkBMHAgtAFzteeXE3A
XJcY8XBG7t4z/rdorBKC40DRTCSD51HRr3Q6PHK0TU+eqJ9ERvjrzJr4VY1AMJpZ4IcEmWyMTXZg
VRj4gastYjkzo2GrnclnhgirtwK7df8Cdjm9xLM3NL+SWT5M4GrWKouwbQUg8Q4O/XMBZT6t69TE
zfC8QACLlyqBREqQ5W04YFUs1ku3qfEsK8+w3k56fjmDyA8MliCKT3Lrmg3R+BtCTIO8oqK8GYSR
Hhv3PmKb947GfWAhqN1EnRVfjbDJ5epIYLEDLNarlELXBZNhKZqUcMqpm5nF8QzWLINpNSNLke81
v2vr+qJ0K7xcwGY7v2KEXvNwsV7Jg7bFBrXkV6Dp7oWccKuwuIH1TXUlhCeWjFx74aLvwF0xDQhI
F+3KeIjgg95oA74RU4qUQ7k1y4atQO4jNBgILMZp0gW29kKL02WS5gZQXapNRJinYI155yAxeQWu
pSNKouIiriiCrNXOaGiZTuuFV4P0lXyKtTizK9JU3unRKGcHz/863I8QZ3bDQZL/2cK0+A92Zaxo
Z49RQDI9LAIt4LX+HeTi93a+h0dHZ2ZCZUf7MX2Fjbxk4vId5VO9aa19Z7ILK6YE9aYgBaHoqt0c
0GFRXBW3Ov2UwCc02SUIQdVMJitF/nkXyhUITsHr9beEpAocRUkf6IybYvZwpR7aytBOlC166Fgw
iot0pcTYhSAoPV9rUFvsmZ8jBuORKCDYmPeisZLPJx7swOOEFC8oWSPNYbHga/0DMYIxxuxl6kaT
4r6UHgRWcoq9YxhY2tcq4muLc0aR4ZmwMD9WwtkQpu/khVgW7FPcYnwEmYU3DmbY7lbfFmaXsMa9
Ax2wYRNZeknN2h2GhgBsgoptFxdceEtZ7XkvFwcdmqgBK3KkH3+VcWfX8vQGrL+5PTLbjFbimXi1
tkHkMFn0A803q7xUEy83ub1dXE54Akm419pVRlsth35H4BIv6qTdRK4BNjjMByfVdIYpdGjehW1v
IPbn7w3DRA2Ye68iPMKzqU+fO4QDy0nC+RVvcKeAJEWAcaHYBNmj2SIht+a0L2ZuLEMEK/ztM7sc
pbhdazhGKpyCMwqhSTSsbrn6ppsUZh+ua/h5QrDPLJkt3d6s5rh32Gt7bRP2A2wqyrC+pOlcvZd0
MK9dylLOpKm8J6tW1dl6P3XpuK2DDtLV4UprXBA6pOeYo+9LWfE/JaEFkBSXjh24CPFp613kYfnZ
O7UdCfRe3NMK1uvGK7yda1gKZ8E2GplDYAGmFjWrlmzsfWW2gyR8P2eFA011dQpOO4ojOlgLp+42
d18FI27FkeIEPza7tC7IELur0up9unVZjNYc5VqdS1XULvz+1PnQNpWE8z97VIynY3OW/UdeaZ93
lxiSWylhok/cbn8RQPAiX+GnJ9EVBM9Bnt5b7qBjaO5T43NzWNfMeNpMXUgVvwUT4YHJRnj+19yx
JCJis0SfsdKXkQz1MRuAvQo7JRYtbZvTu6iORsawvdGudGhcEwckETbY09It4sbwacI+ChK1o0Lx
N4TRrMhAxT7qiV8s4K25dIUg42F1kyJo9zdob36NoPrIewDZCeXe6TE+JGl/M15iMQCm1EBfpx/c
oo/nqv+30iDIwNL21yM22utuoD1BH+5xw33DwsZqjqiABu8DWU31vnM7cbTeqv6Po7SN1SQ3LivA
KlDKGfNvUz250vwwrI9bNzg5tZG/jPhYAIwEYpUW8iIg5GD3N3KnRYl4C6HAuHaDH4DYIn9/fBkB
EqoJuYoHOsrYS/5VYD24YVkPC/g1PShGRX5nGJ9gOIpZCRXjfvC5nKCYnES07EMGrc1AF8wN18qm
u5ZGjKJ1wiMURnhARBxD5TZjZ8lPletRMJ2402W0d5rBXrVQQxJZ/6Q26E4iJGzKws6XwJMOQ6OA
jYr/p3QT4gbwa4HV0AdeHQSBC0Mgg2VVxYusSqHU+kiS+2ktyh8+nFQkzmF4cEHSZ0ptPr0J8n9F
0fSmTQ2jbXPKrn4V2iKJsCzl9mcmyRcs6ZzpGvrk76PU4rdYBtXpbv7KEpz9hZvvoS+fNufug+zt
kheR+8y6CI18uWVkhWL5ULCd/AFsHn9+4a5GWCvPrK2yc3Yt0nmhzL4lCCoP4oWnn13I/KUbzurO
9uyQi52A+qTvKK48tcJwsPYUczyV5P7aMIfBZqfo0OaivKOEJNYdpFxQBHi5XtHlnYtbC9LiJd78
QSwKn0ltcFkiHzAiPj2gqK1TLMTOQshOYgNVhv4d6U5lWrtHMP+DmYP6UxCvRS6bYf3q0zRKYpcW
rlXZa3tM7oZFbyJLb0Rd0h9VgNY7tWMCDQAM+qU122sYGntoEdvGvUtN4gih94anxYKNIMFZWmRO
XsyykBC7wbCYjZV9HJhm9D4c07KQut+i66CSrFi+mS9DSfAJBf/pbGFfMFB7YUNFYMeLXR9LOpfn
aIXAwlUaklJdDDylHJSF4bVwFzPSAgzvc6BS698SU5vZo33y/QWgAtvGKGaJaFjYelsh3BdTRCho
JHmQfcQuOAemNvu6CIJTFWZ9OsKlE66DMW8BEL4cYFeLdrteHBL4bF6IfoyLb60QO0jYH2CxCqH6
G1y3b/1iSn3AMoFEKZ9ZOomijfvvMa/TnZVppDoRk9kGfyx90J3sl8LiDvaN/iCAogqbUsqASlx6
uh3OERwVx/nN99JrnzhV05JjHeU6kODqX0xL+4QGvgNPgYW8qYtM7yGm+WVHzvl7uf6x0sJj7BQf
O/MvZhkkQvffQpxi5szlS/xJvlZWVllGqNm5nHdyQsajkXvXp2B1AZ42WkTYzmUxQAXairiot/+A
44Rmg9Gfym7dXS7WP/uR/EPi901pKG1npd8Lz6YB6RUkosRuC3w79DBjdTuqD9h6FKbXfhjKoRQJ
iUZ8D4orGI6xQYM28hePx4sFPdbZSrdhWNUMsnpwSaL7mL8YBNoliP8AT6z6WykZ5GWnokiaBZXN
f1teXbgZcFOavBnpKd9tnrjY/PjIGYSN97O2cA6SO8zTHYDfWAGNfxQAF1Cu0GMRZHtAzZ5uuZA8
HRys3d/tOPz8zcEFKIvMPGgsDE+ecc4vKo5lLKxE2iXqB7x28adn3owVKA9PpdxneDkVzEMuD4zT
O9pH8tBC7R3PNIb9M97nJ3f7R52BtdhJroh718ipeRVL1vECBvQSKTYIDlkzxuswe4iOmDwgceYb
j4kHsWpbNJiezcZZ55RJUqoDPXsDgj8z3Yln8EdMAezJqXWimbUS3YRSWEz9ntsJZSOeotkHrtP7
5kWOsMOSO0kwOQtIx+RkT4ax/+UlDl1qCubmVn9i0BmiFH0VPjX3c0Dxflx8j3ERYwf/KSR+Aide
FS1Yr76Azfq7L1MMFFyhfV6uYW5aHx0RFvFtrEq0tQcBAWcZDEZ19YdunyK8jcGJExLVcwxfXJ9A
SjEQePLUL1mv1JgiE2YkE1ueFNWHKpDRRdy9FX828gv25UekA6S0CUdEGf5e4vom9QMxGbsDgmvY
cuqZ3MBj6yBsAciueL0o6kYSUnCjcUoLzbjYI2WPQ2QJ7yxUi249EUnB91FS9fMsmJXOM6ZIOyPF
n0/cL0tWwvXe7akQgXr5EqcaBes+/F4Lx3ZlsxHKH8qfe+z1xelOXQBM4Cs+rPlO46974HyzHRcA
mnz7nXMF7Py52aB7EhpeHHnZf6rZyULDoDwn31dAG6/08JC9ydilZscK+aReuS3YmUKTYc9Gy57y
sufZS98yMnCADq96Jku9h+IRHeTJLM0e6QilIUFrANHsq5By9zCJYM5Y9cIndmpwe3uD7TUg1Pyl
8BGqEX55Y34wJRBnWk+PIByEdnnAI0pyqBkUofjdHTWmfF0JRM6OibF6p1royLCja/L+KUsWE2NM
q/uGfiEuzVOoWwSt+G8bPOdoqMnlbSe9GkJEE8jeSc3FKgp6a09VcpwWfyTQJ/wSL/3S3J2QMsaM
HwKUF0BumebAHZ5n3PlcOuA2vONS0OHrQ+BANOExCv1OH+OFxexqVrypVT06SvH17xsRvTDNHt+e
970eVls+7QaWyDhssRgXOnUA4CpbmIAyi4uO1wWx5HZLNQXtwYoc2E9TjUiwlfajhcBw3vLa0PTn
tDtUWvJ+lBskHZFhH8BPi+PqxqLB69ZwD3zB6u3ABuGC3Ds+EJA4FBDs+hp9cal2IBFlDzof9nKd
8uLBnhgklO56uRIPBd7/C8D3bofhhcsrFMnyMjKsllfPsjXGg1TQlvAT3UOdFC+/c9byaGu6Baw+
5535Ec1iGotb6QNMd0WvRUAgpzvqDFjmAo7LZU54q9vy1KOs45AZdJ1a7gT3qsjjrNJBKnpe7pnM
XElTByvSsNKuWZF2hFXHWgrmx7Se4UK5i2cKDPdQ2EEcRAlFPxBLj6Um5r4ghW0xlpleQlpW4YAS
tUEeGElNB7EUKEYkE8lFAATI7oyWsAeHGCgYzVME/CBdb6X+KNDZekCKNWST65k5uoNay+shT1Vz
lOkQ7IsLDrIxWG6nGfXqSdhpRSRLKRFNZMN/lo6ZTuWXuAFz0cMVZVgLY9gJUooljQ7ZsyXago5e
vZfRohJe3hXjj/WzkPTRtzv4sAk/fh/3hQKzZ7RkfD+BwrPbOw5XGNg+5YSvhpvME3KbHjTBCAn7
Q0o1LBHOAOcYGNFJ7PIYtm0gz+BPcECnihE4ISDm0COar5DTxocKkztaO46cVlO9uIvCODTf5SEj
s6ClWabDJ/vXOjAVWJ7RDCB94wwRvXr5GnG8PEaux3afs/B6xC+lLT5qRAHgBu6kMNfKAuiRZH7i
k9WB3JcQtWpvgsy1cL54b4GwmqcJjJqX3I3b8RqEEUgxVN0Qe5Kp2h6ZaTwbyFRKwFOOVEndNKrx
0d2XuWeUMGX7ZQpIovFhwsfUzGxhmTZaXwF8ew3s2nixQOK1PjCv0WejrLPYLk5Nlhna5j9Zgbh0
xevRi8vXUsbzX0PEJyo6yfUKe3FTnnD/Nm2rP+wYtXaCGVzlm6o1Fp5bl0f3uP0I71FnQv2AHE+t
5fU96LY6i9Y5szz39hssQ4hKPu0lpLUCWbF5FySyX/m7xdMbXLDTvhi9Bgwu7XhLr/DawRz5CrB9
it/ot/vsyMNoZE59Q+oVMNJMxpOx0GzYsCg5Uvve97Pm49Rb9vlHYG9jdlotQSfT8IeRtPYwNAfL
H6bvrb0mr1RNFcmtCr1PmngTmS0byWkKStFXkL60R3cszeKGNtTmi5dMq1HtY5WqqHt1C0SePQaE
F7JhyLJl80cC/vbmLvdsEVn0dX3g3jI6pWoBmjHlKllxzR/zESG+J4cRLxthp3kWAPh59fzT36up
PNZAN5yDabj4ev1k8k9/t3mIOSb+3HNejAybxsP85rUN0WDe9RC+7Y+zWwtFHYdDEIU//H4nq0Vr
hVsabNpjb/dMEQ4QUYdrkR9rdw4cjUErif2Gkgtuuv7gygjAk7yrZe940Qa93idXfp1ccm5BQuzH
avdBBrKGCdjLXcPuaIuJzHIKSOw5gTIl2fVYNTvQY2XDpVRBbhNe4cVlkE4fRvMO8ANzHyM8phNP
ml9oOMApqHJ1YByoBPHCFUIPlrJqIeolgqTe/sXAv0A0lM9TtQ++6X8r3kg3htMbiWUjNB11i0Xm
hXfPtwmh0xpqf3LXze5hcbs6+/tyrShzcoUZKMxxM1UIibKafJbQItP+TNCiLCYXmbJzZl152YXY
DME38k0O1nOs+1AQCoMc3I46Spg3j3bXXlYEO27GVG2cGFKd5nifCw24HUN/dcLhAigvnRrp8T2w
hw9iqkEIy1J2TM5TMRQ9dS9NaSwTmGdPnG6rMK4A/ZAot8fJpmhPHL+dvZ64gI1sipZ+KuhzC8Bh
2bB5yA4EGtrOhesPwDDOTUdgu9qOz4uSgG04DepthSh0gY3qhufBK51IE1CgYtLJOaukJVOWGVaK
ecz2aiJltyNYoyHutMwIv6i4iROXUN76x4h+TqJAHMzbmW3ifgoB/4pOpTL9pLyLH0T21Ih/Om4t
AJLOKqLUWHD8Xh8L7BwYW7RDfd3+AnEQjKiJ1ZUHbLZtxFhduyL/myUIgxAm67jkThixotYNTyO0
AO1KUFBPRzGhTDc69Aa7iPhvQOBRr7xWIPL4zHL+EkfEgFVHq9H1WAraicPdZFvQhwzCpC9E88Ab
X1dA6J1GnPjEh8kH69ZHzLc4z8bDsiVyc3EUMozjWDkT0bPl0/BtqFvGloeT4LAUYW5JzsLUCE7G
zlKYacuHjCXmDjmXYFeTrqob6ZsAhe/ScJW4xxFWs9A4igtycqvQTzymlmrtihFguxQayxXTgT6z
GOxbsmz12h1pMJRLalm9lWlT+J3FWVD5/LoGmdtdmYt2T/mqyLgaB6gLXDuWd3th+EKyuBjYUvvK
PmS4MfFlXtxZgnRRNeVcY08OdTgvdjRQAsvc4jOCfBs4PqjYYqETcL76x64IPTcwTRnyfwWwn4g0
emqN6XwkT6shLF4FvqK81JeEn398FPs8xasWiuGBD8EXUDsL2LagyIzKe1l+EMhzDDrO9zWl6B+W
7iuB1671CJHUiDTIfbbg4ldoRl5dBLZW0iVd3ebbQbBbKXE8SK5iLOL4oi6nHxqxWIVGvqLgOYvV
fXI7mqpSQHDQPcD9wEnBfqSP3lEJUK+0FT4B0/2ERFdsBtiythA5EGYsTu7JkDbcqwRxdaBsVnUr
BpKg1HsSG0ayOHroQmgRbgPFN9bHkM0MuV4LC/dkWt1vrFNmKkSxqWNB0Hsm5+s1MyP5OPw160fz
xA9QVy8B9hQwFpzOeQfa8r2hPKbKilmiB8YIF6fEHFCgjZPL5WwpnzwTZ0wOp6YxftT1iy0HNe4w
CWXLQAyen8SuGTkv1aerwqkXLd//iUCwFWyQY9szLwCZg457ANfSC7XL8lG/ECgCZM+NzjrfNDti
f4Q1TtaSNNhku9fw04cAjKBIMx9zy7wzrzBidiWEEJ+9V9hz7VEy6DWL7e6yYT6ywiXkT6tHyZnW
xV3d6+vwKr6nGLcfo6ez/cwH0nFdMqwe+3iygvdS8Zg31AH4aQa3m3TBSbaRLLgB8UI21UDCFxcS
simG4TcRwSeBWByVMvbY5eGEo38WMe3SqWu1rqG654508iDbLw3D8sFzzD7ubM6DN1lPeSmcd9ah
GWT17r+rhimNdrvyYJ0oPhuN5JDQzVnTHqpMMxL0ezSAsxcBuyPboNmmAgneAHvX3mhaCR7YLuNJ
T7AwsrCtuPEMrTmqoe4JscSjyHbMY/3yp7nojtF/C/tW8q/Hn4PN34IroGnc7jlWoJOus0gLFr3I
uJROgeTd6BKvcaZPLAnFD96u6NoXwTA7LNjuwNiiuy2UGf/BBP+rxwBjWSi/x77LjAiFlqAKzT0b
5JzNH5W4o83zAGsPnSQPm1m18jbh00gOw95AdfCTj6p1i63Rjs/+oEuJRJ3aY71BTlmyrDI8pxT/
fAm2/v7IC2i9yRjLZkx7yyjzjbNA2TN9Dvn+/h5ASlu0RHqOXgH0B0VfSm3l7IzkKZM80tnCcnA7
218Wh4b89spTdk2WruKuAw9QVAlexmpU+Sk9TijcK6hv1KZztopz7jFhNQ6rdIpdNBE5Di6lCPFx
38dO5TmefQZfPRtObUoKXJt5N4Sz0F9VVp/hP24gXrDgQJueP7pJ/RnVYKKpX8i8SnEO2LA88WXp
39IpMdb9zwIBzdjvDvhqVzt2YOkT6jAgy/1RkELhMEsgED8ts1Za3rpR1cc01etYtu4doyTelJp+
GD7cOs16O2sKYkamNkbjyKg18il/jCs575uIrWvTtjoYbNJsf63mnTFqoVfxwcw0/9UUKKqBRThf
n+zBykRDLKclOQ1MlrMsx8iKXsGKn2e2lFgeoEt3J00dFoOJAhAFoG28f27uvhUqhYhaSslyZGCs
3zyKONbMlFhjtpRvSC5UHNHu3wNCjyJdqjvwLngtFdOEdKgjCrJQaRG1+8VvNgrrbuHWbh8xAwm2
Br3skKqzSeOMj9YOiT2E4XlXh+J3kykQLPFi6TkfHggfCOUXVMOeVYcx92GRWPaE66vUV3EmCd8H
HGP6Mrfr0473NcXIyaKZllwj6zFSqK5r1I2X0wrcSTrl4ZKfC3IFGSka8OsyA+f/UhvyIA4e2XMD
sn7OgGoElEP1BayYKu6WX7fIpnt31nUwJ8IRP0Lag1bj8QGWd5ZUUbH64XCZtGXsPSVW0cG3rkGN
0LjESrRaSdrBkNkYFiu2wOa8sPhe1gUoHnP/RBU3Y9OfNqnlnyWMLdIPRMMCjTVXkEnSS7hoUx+y
a0i9rcz54cKTiyg1Cr15nY5a38QLkMliaM7w5yMzVF3N7KYQUnK63H/DYI5jdqyfQoou598n9bI7
RfyXd2mWewteBX5xGNLiAq7oURprDm336+2NzwVNDZmgVMGF7iVZHC8x+4ed0AU9/ZS+31r66oyX
zPr7wD6NfwFLAOSg/qFwJ6Ch6rB98YSDErNmmFNf9LtIIaXStT6FlC95tWieP9LPUPWT+jn2ryJZ
JvFBMcYrX1eeg+B+Ajlfr1bAFfpMRCiFP/EXIch3bP/j0MHmtWqprPJ0fTwGb60Jqv5VBBShRONA
YKhqLNSwkZuWzyRPxDGCzOoJc1wMo9t1FJWnuRI7ge/N5LA92E4fDGKEY3fLC82oxg6zdizovdWu
1cRFVaYp4t2Il2Slz+qm0ZFtyiwQQTws83Iv+ZUEjbke7bbx4axl/tBL0aWp5cATpYNpBvb18n0R
q6OrU4wYW9D+jHQEWvSTC7V3iAvmcVD3vWf88kgpc87pXMoT3Gflzsp1t3AuGUw296bRWYXK3iAw
m9X2YGjSlfnESJfAbpLYGMVeOCeNd9BbdG9yXb9XNC4E6YmgzItrTefQsLJTrkNa3u4GzfBAL1rL
15Y+Rd0xGJgI2Tocbf6GlnfSWE8lssHfiVzd4Ka+nDELKCGLylnvz70bAHJc9/0wjFM7zEksSoC6
F7OYZ4Xltk7MGuGT80WgNCBXUtZ+Ly0uJbcPaeNbxPtbS59St81AYVC5MERL1llzDsMF5d7r9vFU
lnKp16HPqSar26WiZiLK4Aa2MG32j2IMLxfVsSY/BwL/QMlTkL+J06X461/pLMMSuuz8yFJUdwzc
/HDqMDDl37VidlZAombjxITPu3veoQA2PTI9BLx3xiax+cNV+FN/uc52afhXh4FZg/scozE/S+qi
47PP9ZaxyHL0tfNbWHPwM985OVaikmUmP+xpFkHyK2HVLlOYdV9pzaaJlJ7a+jxgbv9Vv6HtCqzn
LyxCQKYbT7xl9EULOwL0MppU6ILo4fBnZlW19JbwWkNVmrsQH0x9PZMPkEqb4vvT3cFeDmBjK65k
KzPewI7nm6NxkA01e7YvbUYNjRBD+4ig1ye6K50DkjLqBxZbXLwaL+VgXQtJopgK8i1rJWijoGVh
xCWaXHjLiKz5gNv99jAShmyo6GZfxzioBpxZEP9NC90Fq+OkK8CPUFRIaYPZz5I0GXcEp0fnYJY+
82J75sjlGv0jCFOGEbCr5FGe65rNWrImRRJt0QOu0udmwIWbsvEEGrsHKk+aKk1eJqtcn0IWw7gM
sGzrYJ2YVYMtxNJ/0m43UgIhdI7K50lVU3O1ZKC58o9wBI6n4N7rVsPpcWWp+F8xbf4xlWQtJRj3
VNrzenmgvAFPv5+L84edhEAllhGJfj5gczC476eE5ri1YxKQmXa0YP3+JjXL8720q2/YhXTJDfcT
9Wf4gbBj5x+8qRrKVDPyH4fUZZlFjQV1D8dnL4BPhpFTVA/XY0cP+1etq4f2AmLrq2hV6GpZaQEA
Vd0t6j7/3qUClTe03oWvesN8QP632WNbWVdkAU3dIAxlDpmfXxCJ+06KI/9TTsHUeIixc6vh0nxX
hA04NKOEHxFmrtRnfj8GEh7ppFDHX84evRI0QWOqIC5BobfUw+QZNofBpeJLjsgfJfWNPRNjOnEN
+Ka7NPfmgGDb1ODpjp9vRwWk5eK5Ne/GrSGdSaRHTOXHORY9j1VS4EJfoRFcKkIW3FSigQ+Dv5JS
2q1MaOlu6mGE7ibb0TjbSErmTmaEV/OPcEdeE4nvMqfoMiL50KrEPo6E/3t7eEkJ6vZlnrUJCj1b
dvpPkC9bUB43ftk/YgpBUZmcCI4uzc4bF1fk6MSdjdBm1jTFthb6Zm2BjrRpqQuAAduOo1Z8Fq4s
Cn03fYIytJE2F9g1nfXc8zPKWJgeeiCdRQKrjTh8zzbfOCwIOfbzXLF/cMqof+j2Bq6FtNyHRY3Q
HrzIbXU5vX73HV9YfMi7Wd6o2EYEem92PsuuiVLNzS2I4qpk1PWeTJBHp+zAV2vOwZ3RY7YLwBgD
xEBjoRDWjRPXq+xOJZBk28vDdisBNMACPV/tSSjsdTVU41E/i+qG/v7JeDd8gEZ5cQdvkc1Pdz1C
k0fwOej5Xyg5EwQ75qD0vcy/cadUgOOa6LEJtyjhVhbnnRJxVUHgh9u4ODY574EsyxrGW9HaAybF
TNlYlzrZaTVVia9zgTtpW5UtPBw/1aw0J1pFkIX4WmT/99DXB2xEDNRDr0p7meBTlpDt5bGfZtxp
qX8tErrpETQ5FXWsle6QsNmCx2KQ68Bbt/In+OrlaAryy03w3Kt4kL2Ar5Qj3BDYFSIwYwwIWfmB
l3CdYRDm10igI5BeFwIYaL2KAO1wghFNVHSm5+hSyJP9TLzSgiwS4LMwV86YAAmXSyMI6kjUzHV5
ZQPABPoSu9r9KGxNyNhuB5r5CBhGttKAbvJKCFnxqIjTvbuPjr1vrK/cbJlRt1YwDhK2ezjtlEnf
pbFg6nuQ9Ncy5+qFfehUQb8PvWcEs16EAfEixXWXo+RCRix6vJEJgU31vbC5fmbrl3WtMO3NlY4H
t5qBT4CKnuzAXEJNQahNTmh4fphlhfbLZGWRz3vBd7QaUgOpQC4CeAWBxJarfRlOmZfI3JXa1cB0
XAjXHJO0tcRmj/lTOXSwOo7q9faUBLJsEM9AOyNSw+6YDVjuA+t9nYxgED9k1SDdyOEfMNmpN06l
6C8YIneChMHLF6I+EC0A0uvAIeT46zYXH+//ygDgU9OWJAu+HEXx7yNPBX7tzxkIJqKSboLnqCoK
wHO8QqAHP68ghJ2G9GkhdjrLqtlkTyyOW9unr2o0uSNqVCnb09wSiRzCvCb2irosULP7D/r1G1gj
56xifUiJFnG7dMNv1Pev9JfqUxtTRS13OoOursL18AqOzSeEoU5W5izWDa7d8mnkpX4fvjWisYpc
MrLR8x+WdxvEgoexU63Z5pZ6gVa7/Ut4HJldqj0YIDs7CyHCwDG7xH1wYsqVb0iAbs/Y7r4/yn+O
IaAAhtOAr5mhTWZj1VDiUXk3fUC1U6HCbdFXts2l8eMtSLk1KGN7FThDAjNAKlc+G9emNmczlfn4
kyekeXFp9JT1ZRkeVDLBeM+8RCGKrW/DPYBx86e4oRcNc1PftEPeEFTsvDjYe5zxefSiEgP7mBWx
UDFanExq0CO61JHONefI2GfbeNiodHMn4ucrzrJH5QADQfn7/DBB2Nm6oIYh6HyGUXIIUqg8fR5T
TzJ3TBm0Q23nEOIutKSRUXWqI/TG2bN/UHEgmLR+tuusoZdIpTO5P3QPbzA+I3GXHaYqCmv/Wu8C
fY5wrCNjUB6TOcGqGmq0Z/4UFDUZ7cATG4WPhFrkSBiO79PdUEUfaFyxBZxQPJcxSAlg12yAp7bD
nb1kSbgXn3K6FyzgletuPpw1ACBYB0eiP7xCTXZ0kXYDlRi5gzieeBw9ONcabFmor8r1xuCynkgH
CyK5WwswvdDvzvmNzd2OvCJa27albTpSLebpbvc3nYJ9mZL4DUElYfmnv6DRHH31bKW6PPDYLtjr
+VIg9Ld7hwCVj9h0djuvdzJzQMPR7qepK4Q3XorUaJJZoqMM4zZpGZqQCHo4Q4hfKypji6hYd5y2
e9rMozO8VqgBSxY7HdtFx70YamOmwK68wNmhgMLPs0/z6gKuuHd3+G1PhuAQ/Ry2aqekYlGZzb0a
ghkNa2bx2UHy7Dv0FUj37SDvm9YkUgF5pw/Dr/Ix2IepQxBeLRYEJtjFVwVjPcDJtboOaOX7L9Ks
hYXzjXB5xjZfkNXBXPzDRtR9Zu28OZPNk29cKxPlbbsUR/sgTuXFEGhkrOqwVlQJ8aK3JwNpQszq
2im9OIXuzvIcbqpeBZDb+y6d5T8L1ajORaA/4IrnunpeTSHbGYKKs6gC+lxaj+u1HgPuxN3vUqKO
G00mN6zSF0NEmsayjtp+QM1EPFneuzd5Zp/lqtdCFdQKB2YZ6ESa9ai1Lpb4tn5NA/ahWh5kPDgy
hRmPSZaOKo8ovrDCQ44/C7zRUBOVSfVcgzFrUNMZ0iPqAE5J+cU/GjpgPJ0Ao65haaJaOojILHp6
ZCVVK7Jhx1VxeNNLNdz8GkC/CjGJiSvFeLd1aIVPJU5gRuJr38shkCcKe9jIutWIQ/BwM/fVWYXE
vctJTUP+xSjOJ5VjaxYP4gXbg6x9G1eAo9kW3xGfGozQDRyvNAQNlbnbUQDJ9LwErXeOq1h2lw/Y
YX/0M8RZIGH8nQywS1MFUHZXK0lDdCzmYUGMqWXX5aH4wDigYaETBukEEqv/ZavmlKc/TiBS19ls
Drh5Njd5illBS071wFruaJ9A+pHKwqAnNfpF6ouC8F2LKtaFTQ3uMST0dx81qEnHqu7v3BpVrxZg
hTgsm5IV2pMb+65yqTP0eAIZWp253mRV8CPlCMwdrH9hEjSCoDTQPcTfE8/Z5vhsBIb1NADJI3zU
UwBDxPmopdewA1kn9rGzb5m1maPuV23qqrihKKVH4BRgdTw6UI9QAD7mXg0T1Z6wsi86Jochyr2O
AVMQ8oDEkWRwnWrbeZTOT2dKnJRWnSJ7CxREEVBo8ZqlrTwMGYuPbkaqIFYEx7M9lkd6upTXnPOB
652+BPfxTu6D8KBroYhB5qdQkDFBuOJM8oKBx/GKHrLVrKGpm/JRiF90ZVxKl5GF/oIo/+8ewRk3
KRaj4lVU0mQc7D7rpAYtOOquXnOWC86QpjjN7mk4OPrtGTVrTPIHPVT1q/0H0fvqtQkZHgExzh2V
QtdPd+/hof6+gQX++jaWE/lIivvi7RPoU54XI9WupQOPuqjN3SaqSv9Rg0xQ065n5EEElGmfGPZt
yF5rzZN3egFogGPoRjgBAEbuECK9LGGlhgyMBafSpkzJOiyXuppQi1cp2fmKcSPR1inBaK0Hi9ep
b1VzH3AlieIn3tKFhyueCUc3L4Capx8msvzAUnSRndPiv9XoDDj2oSAaTnBdmvVs/8DhQPGBleIx
rdLU1Bxzcsg7omNlAgA883hqr/OhYuf9t/6PZK68B9zrHBuyKCdqV4oOW/JoELKHDnkNI3DJp5sg
/u25NhheWbKDvggSD5uqdYXTgnkY0s7YPd6qMJr7tyXwV5URvwT4VEIToNACVWjvU9jfjbeSW1Eb
CaBS/Nwor2Um1WEJQwHGDnYYkXnannABmOBi4bdu0lwXDJ86n4vJ8+jUcJK1AubnWO2VdfsOFv18
JjMvy3Zg/1aiAOAUa9KoEn/qIDjMmAy6CCFE9eUOgfYY0fm9srNUxoIkbjXTvL6YvI2dn2NCU1cy
eer2IuN3cnAO2YbK1w6IBeIZDqL8JfX2cKPIhOwEDxgpvQJ6Dpid3N0mRP+0e1fGV1auPdizDmcd
Z22v/9eGsVb7fyn300MQfvkhp3jPEuY3cMNbZvM6Cx9Q+1aRQSDKlc54vw3kXiBic3rboF/Ml4sU
skTWEPSpnUhXM3YKABx75utho54W6PjZl8VFsr4qWxSj/elZScDOzyI0+xIUTC3enfzY5rQ6Jzeh
h5FD6OFr4WcoZgabZIDqPGwpDhx66yammHcnLfhSlH5YzhqhGyYHZjsWVY7QQgEWlBRTmDIdck62
CWEd4/4Ld9ikOrOLYiFAjKkJjvaa/dVkUa+McMYKkn0EKoF9hB+3cfPLk6vT7cP4T+m8aeFcpmJQ
UJS/oPae2nEv6Z5eJgVcwJL7eYkS6Ma4zMOZ+stZ9NX+zSwZAIUmNFBeP56S2cTddWrBCrLyT2AR
so5qhovxeZImHtCT+QLY6Z7JoeZl1sYyyTtHJV1NMduAnh/kl1+C9JAgRm0+0KqtHcqF3f11VC42
MKhMCO2bHhMG+8ES36i3uCNELq7l3cssmftYJYw0lXLGk3P1ewHvaO6XkV7OaaNjE6H6J8pCm9OZ
LNGrFmx6BellZkBSEyZ2MqlTZmCyL5Jho7e6KuTBRMe69obV4yLh3OzWX+Y9nV9pAb9LpsA1CbSK
IAKGfIJ94FmvwAzpUh5wlN7ZEraLpQJf/I/mteR65YGzHp+QdgGQ9+wUR/pl2vGiGDRRF0mrGwgR
gOcaKSG87yPujYrPatJZ4k4Pa+27b56N0iJPrNx/hUdH2uoVgFuB4mgnYaeCa92yrYNQ10MaCQrV
HH67bWzFU9aLLZpxTsJZHUraJ0+IDNp9uWJmWz2+8MhrkBrjqt0KoZmoNYAiMhUMT1vJkXhwIHdh
+4ScT2/lIU2xuJ3EkCYo+wnRteGdVgWXzqrl+CcxLdOGRLYQNh4kvv+GZwVs2cas0pG/zwM6ZSBl
H96q27Bz9xLwhJS1+jTtaXyhR1wfDymwRnrY6BIAiH4W2vO+u83u9KiH1LBKsDf9rvey+MJhdIVI
NkeHYaeKBWYAjTdpJwpisKFqIa12tsJqDlNasi62JdkqDwT1t8tNY1kblVgRGW93NGtqU5rJrbxO
jwQJ3ZjMagvCpMdedfzw40s9NdaqbHcg0rAt+ZiF+R3hPbrVIQ1H1iw2ZGyllcdLlmdjb86Z1AoP
xMewmKuSlAcp+ZsD03aOfYZtdjqnVnrVRS+8g/pHTDZWOTQ61iYO0YnpKNJZdMaRCAvjqbAzs8Ly
R30DmjPxFgUePF9QecOnU5dv5PKh/B1TpaEiJK4V6WIrX+jSWZTnpMi17gCvLNXxJe+Rvmgv/1UO
IhMqlUCuCvtph0q0uB5iuWebW8lOlXq46S/tJgHzalK9U02f5bYhs2e3/9zLeUsJ4sigdvHWVTaZ
OaY7s0Iry5FXUnwJeOfok3fHFAXxDDcX2p5H+sTvScFP3JaLJkxdXPbUA5bFUlxeHKSiB6yNvsyU
a19fK6oos8dDSS6XdPk5Fip/6gE+VLGnJBG3TlegcjkvGxzMjYlAchaSU+CqdtZYNDUhFThhIW8F
IgmhG/WUIPxSm7t9C18SS7X0nXiHt+PFwxy7EYn9/7PZbINosg34IKN2Yt2TOBvZgzSN2CrV4t1f
Hq4zPAcCGjgtgNjbog8EtU14U3v5NxSj/S8buBy/jami7UTun+7YJqr/59v6BVb2uU6dR4YANi9s
yY2MhLBqC2CMK2x0ig8KfoXYs709K2lJ5bvz7p0xKEFtqfSqQyK+dyqKGrfMlnlQMXMoIniyKV3v
3VVu8plTWCqFzMZGc1zAZ5HXC7IseLg9Bs1fijeVRSm2JNIKG8A0gfKz/nzmMxx63eF+BeiDnR9L
8wuc+dW2fjeIdBskERbMBcuFuo4y6V9cqrFDt7UTLJNIol6opvuj/H286X/iwwDfN/GPlMlmXnL3
FYlEXQx8uuHKSGYWj+ZExXzz2liY5GkbU96WM8OJ1ZLfnRF0A0vkTkdoGvFlcgy9QHNwNblegUgu
f5F94Z2kovgIA0um8JJ/A+ZPQf/8SVYkqR7XsF77fSRVsDZpceIur2XACl2ZbPU+nCpHMdg8BOGe
XvcbeRplBGrAkJK9hq9XBjInNrJMGHJKT452MpvXl6XpcdvT11JEVF1ku6K7Yp+FPgnj15UVVAuq
T9edloKcyTbgR8B7WAy5mG2Bg6GcD/YFxzLF7J/AC+Ejl/QHgMOXd3TxzVLtZ5obI1+80bqEIeY5
1cGWfTiJKM+AP/lx6slYn7gaGbN9G50i5onLRl0HM2eOVRxIndOAE3nNqbwM4VTWaVS9r7vk8XCL
e2WklYRQN6FIdiYZxOh8oW7M178aoKsI5bPrT96OEKzJ+AMNeqUwCQEqRfsIyxPkP9Xwumw4riCV
Vj/7GMK8Y1Uzix0lOSttZoZ3hRzrpJ2yGp4n7I4UMLy8l24DOcX6q0tPEBCgtg/XLW5rR6C2tbwE
cFi44RjLdF508Ko5vP1WIWAHrDZq79057VUtorXgFbhtaZR8XoZKmwf/Hz1sl9HCCOJZ1aKP6r/t
WdKi4y16WqxAKQWHqfq+6McTROm3BXOVjccG55Ag5UiboPTygn5ziD2dXSnH697ME4sN2jkX6FTi
N42ALZo0WNwXRUYzQa1WaoqLKYLbflPsC+aqOAA0rLoUBuJriOTVzBekHBUGVxpJxMjqnI/jDkgu
mnQ+XSLp2BZ4Z9A8HpzsM57mNFIKeiewbRDkB3Ue/SoawzbzCdyTxZ1sjgV9vDfBxKnnAzWwgoMK
AhplWUAPl2AyU3FzQMCZqCCUl2Ho54uzwpK9XUJ+YyKlkDJUA6TSQkz+JtP/rl3L5H43qWdVYxYp
h3qK7A77IzC1/nhHj4Rpa2L0CkSqzhpFrJsgvIi+RtxuCFEEozsGU9YczlyyQI0PA1mh91vEjZZq
M8VOQnx0gVocmdE+WRpcpr+7LnUJQ9dtxklN1zfCe/njqcIOMda23GUWGN3qt7xGB8iuLTaRyEcj
jHq+8hClefDrjMWypyi+bhyVGjGj5nldnF7rkxLRiiSb81sFfIBICtDNqnQZp4EIBLY5VvTP1GkP
dEULYhur/oBIK639Hw6OuL2fPyxcINbXwpmIzx83iuGMFtkYSzhuvIEGWKKy6CucYglgw+SidDcH
kA49ScdopHwZkBuV8xUmAdqx31ZLy23XYWfTczqGgkTofFivaFLMwEVnFtbvKFxZ8SNN+2IrlEQ4
TolaIc5B8xAiH3uABzf90W29ybrc2zyUTl7zykNXrceJv2y1Xsk53bOufPvg5ErUdPV9GunzYM5M
aRv4mJ74Zh0OneJ9Hvd7ql8YpwlqxvRiVTFJw2ULJRfcJJyhRSJAxX5Q0BmfIjhLyOE5hllm22ks
GmMF/CG+l2slNeDaw2isef+cItzcK0jbNoeDteKnIU9494oQaFH4lq/OEivDyqPPeH9ezjTDqmoa
qLcPhMzSg1XNzVUMGXomw/XQDOosKfY4fcD4poKFO0ckTyONMIQrj10wys+OqWlzXTGJ2dbYoGmW
fooW+4UAv59M9UzHg008wO61HTVBwy6v7xkycwgmElzfZIaQcjjMqLbr91+kunVJ3s6TAMT1qC7r
GmKlStMaBzrbASBmFmwljF2Z/Ets62coTwcauLycEdDn1tavHslKbGIKPrCdgsNvqSc1BGQb+Bw3
1Lbvx2WIaZs9pXVA2A0KzpYwh+PHk2PQkzRwA3LiNB3mqKYoIIWpDrHM9gw+Qr6XrYcdgr/ehKdi
2I7Rxt43i47WB7SxtZ1cvEmTRY+AOW+x2Vzz4vX9ov0ugUiHsUoD5ChIFJQ67nOZUAMAmRlI4o1G
kX7+NujVcDVIEnr8Vf/HcDVYooWLb2Xjygo/g/8yLE1rNsfYJz6mm2SwtuLqWpDr5Els0Wl3xFzf
+dODYcfSpEfDF0mDGsJNhUkETtRFZMEgZakCmThxltzkVu8a8JvoPgTKprXOFMTJuq9POFad8rKZ
dxKMz57rm5bGKdDYLprj5YoSDdO6caQvMiT/z2+djz2Y++w7qf5Wo39D2CQ8iN8n9OtIJWYIhyB4
P43h9dGTOY034YULfAZIhmmieklx0EtnGB2gRM7zI5BQTjmEAOO7AfqN0QXledaFjeSbSQlB/G7O
0ie8Mll3NVrmGnBydHOXPh1ZdOdYcTxDozS9mVYHYQbJ6TstQVfK2IiJdVnVwp+cJPJMxbeFDVTB
Abp9/XPArNGgyYbRgplXX5mP1imdcScVc2OKm7pIcEPURhcHnxphVf1BjrwQxeFS/ufRjk+ttH9+
dlgYSRVGnFTiMBu9XTMwnDBzJNMg6I7gr4uBt+TMd9POezq4Hzc/jgWKUMOFq0KPmW46FhWER8Op
FrADKzcGipdSnjxE00KTTbJv0ZWnZWhmJ3Dp9XIMmrCH7cGfVS3MqOSM8J/paW53ayLjRecIp6ZR
qTmCRJSwg0uCY23a9W1Vhht9/qd8mOQkqZ4aL8R9mLjomHaQO6KcoTJYPOJSqxWvscwmAToIsx6p
Anv2vG7rGi5fnuIFonvkAngDQbxTIznXBSR78QVo0O3AUTTOCOZyb2oOvtiKD+6I+2B1TphP54FM
gZDvK4yC34bzplDeNWVhqIu1Dbbqbgq1+bsAvzYHTcoFk/v6Iiq4YnLevCf1cdzudu2XqV3ysblS
y0j9hj1drpflNZcNP5LOWnJL38hPSktS2Hd9NHzhOh83wixVsjm2P7LUIjNUIRmQwVYdZGRmDFNL
BI4Bay/9m8Nx9JSUqYKB2In89Uc7AgsACMHAJ34ywM+SnLsOj3FoAUzF1YmR+FoSloaggykQcoCu
cq+VAeKKBDVjAfcyLbH1TH/dbO64Z03/ewXO4cT0VTxn2mOUXKISLxho0IVpGSYheKlb1nITTOX7
C/TdGFP5+Yc/MTbMLj/W61wtrueVXq8fdKlXmSjQHuUH5EvcdPTr3X0btjpo9YAMa0L9FwVJGfuP
KslMTTULadqoHWhfsjhEh57zui7Gl9uQXWm7I6fhWJ7Lwa7h0n0A5NquI4q1a/3I7yAQI/j3t8SM
O14/VEML7ZpUwlRFJAjTqZgRplzbkAUaauhljXE6V4PrXLBvKNnIS5XUiS+vafrPUX9Z4D7thIkR
Ddy0OVIA0yusyfmmMQC8s6VKfVAcVhNztRzgpHgQS2snJMkX+lV6Or/opKmhBs0RsJ0CU+rpjUg6
FMFBth1sTCucAAz+bRZ+0UTPUtFSSZenOWrttYZ/JDzFPjHbeUWzDEl00DuDv3ib0uU5PG/r2Sju
CSjn2gEWCepYa4TtZxRBxHGrpibb3AZ/h3G40RBHN5VMYlxs9pPzizKS99wmVCsJdgkmNnaCdyNo
JwMxRIhQXz00vaxNGtzDraWzQ804xXbaiPIclrGJK3Y7G3Xw042we6oSCwX4IdlkHPR9mVflGMsW
QYAe3MF4KyuIkwyKYe1wn/OoAaHrORrP+sFIDO4T3QL0O80SA8NicLCBJT0ImUg87kKpFfrDSoJ3
Z6YyAB8fU0ZJJrQ3f3M1FScs/ZE7Jppa9+C9Psm3mVMi5le8jaw/e7POQjcVNQJhslGKBdXZHqX4
f1bAy7zmhB/u6MGCTHH5tsh7a8Q2348wJKko5DyRaIx9Z2qfKriyThOq6vGGGpGgVLoIOcJkxnll
dDgOK9+OzQR2GOyxn2Dn/3SOsIthofMzyoZVVXQOlyx+6+P3YrJGyIRHgW6kdcReV74BbpcJrgEO
7gUq+H10D0uNLN1psySHZ6zOgfsZZf+19NJlwnTWcPYFY60JGg6vnwXtDTrTWUm8z8V3VuzxlqpM
5+i95Y6TlkZJKDA2U+CJuM4/HDuFiZSqFHkj15fH7aP0TA1HpyJelAg4DHrwiX4Mdy052s0QTx2r
mjskXDeiZI6DKEiupm7nbcl5wt/M9gxF09gVSwJkQxn0pL/xJFAQVPxmAzws9CVyuE0XZUECP3d3
jceZaKrmPyMqF5cbTQcls0YPu+hjYPHXBUXE3Gc+7IQa6lXM3to23E+EYo0BZSX4EcmozDheq+X8
N9D2GnALFsGyDmhYQD68SDh/X2vBy4eUK5DPqiR+ciotJWiiSqVfzYyjZkaeYpPqn3+rdQMWQogc
0JFpzno/cMZdRDgt0gfzjbpvamgqd+bKXkNfZW3klm/9CbJA28r9up72JglOGNGPnzNj1EvYcYBP
5MrJPeA//B6Q047dNcrunVWMZ56+oCheXhiL0iBglcaD/fGEpwvfVNzmwQkykvg0lnbkY+2IQp7i
rwPLfcXqJUAalA7S2rZDG3wJO4PMaVjh6bvae/c6y/MID+vcdaZYr5Zc6fnjL5bOaPv453LHrrks
Zt3MNhEz5QVZCKkS80Z/l1vxU4kO9pLqNhmfshNGsyN7qQYt/JbiY8NeulvXDXOy7Byh8YSlsQv9
eB8vzxJB+6+KFndlnjM9WxNp7Bhr0hS6VRjyw9ASOb6VlZpKf7qNHcovmeHxabsdf7eNHrHk7OOg
ymi1BKrNwLOeM3KjGNJnfbw8Aadaf8bzYIF7JqA2NEe65JFvfu+xYXDU+Eg+IBwGKRNVnFYy8IIh
O1P4n+xSN4X/DPf1BXj7QgiVZNkHCctlOQoGnef877FOix3hLc4br4YyB1b3Gz8WTD8pXTTTO1eJ
B4PgrlNtlb3HbCOe2GIKLKBE3rPMGHwcRXjQXMDUILUzomIJ7sHIbR+vhJbcEnjE/FsbcEN9P6zG
K0DDYY0E5pcZiqqKEl0Bon+dbVrXYrsaz6CNIYnuNsmrn/1Kf5wpqhd+SA2ss1fNId0CD3RKKJ6e
hemSs8hddZv66dBxMraFR2dND1RCfrXtIj3ENQ6AirzV/ejSbBK1fyGGSZuDyhV1zsUlFZHebsQS
pLvcSyB0VRySxKGU1hPptnHPpARNBmFyE8CYCwkvAh28/5GvEBOl6ahqza+ohBeaHInALjVouvaK
6bqstnhvxyRrS7dVCHrqZdSicaOIZfkQRiI6uhfK72Mspi9yLRJvP0BetTZ9mEgBCYwXud1FMIl2
qWy5I7NXnkO2MX7G7F3o5B+CTn6LBgqLm1ujIFoyoeF7EAanR8uTwOVRnZosQJCI+VuDivTEbqhX
kyAhVdU2BazcjrSM9kJWyKUNCDG2OBHq7zD/lunCw4+KfB3IzrapfqFFXoKwQtcyxxMf+97w2KVf
3+JHnAByx7OATy8Kyt0L/3Ew0rdfsUJghNIRYpPlR5Gm5cXfHwOEMOGp9DrxFlgz6ygtgy6orYOO
GnQyIn1owV/TMDMUNGfesNQzuo4bZU+7VtyUFy3dy0KP9Bt5yWEMIDq8Gt0kUpH//yRpm+FMI8Qm
vdlJP7Q8qZWPDGYJrLb2o573rMlAHAGyb6Lgo3Ev88CvdYN9oiIfnmpDvEJeYmFCmQAevFjtWuCz
UXZpJfJyQR0NH2s09Y8Gg1VWb2Pv9N38CaPGbIjfgH8ad0sIySKkPJhRuc8kiBPU7jQWjIlNajDG
2hjGcBTsHrNhAHZb7eIhC1PPDGnFxrky5SCJb5OzCk0q4Z8R1FCAFAFKYSoXudCjxoExFTYHljuh
wCieSB5yLZD2YwE9QwDiNY470xCzzWX96YP2KuCb6Y1Ldibuw0oNzktrJHgH+U/a0QT57V1i/viF
Lg1+M+Cd+9l1CAqT3iygjG5uGOzr1p3Ao4LRi8NssycuINCQtxYxihwa/ZP08Y26lj3qKvVjNTj8
SYZaHqrPh71yvu8QaC9X1WOFPyzlLye6jCxGPQjbSiva82rAq5BwRBJYyYh2Duy1OpJxQwTfp3en
6HLGHx0AMKtPleGbQA4eXlVpy6vELvzAE14qGKKzMHXTwYLbr3StpSIKr0HsgBS7qpZhY7lWkdlD
ToF52AXololLyWLpJMatzbe6WNU/JuYO8OQL6yUIjnJa+054/lqRLM0RkdV7JJnylDDkT++Zws/R
ZmCTIhbEunOTNqfHx2+5SGYxq1TJSKb8Kf/htyoW/l5FaXXOZOZnUZI+i3qlbZpjl+GteNx9P/jr
1kw8D+Z4k/TYBaGPVOepvUij1bZRxoX9UZNaWXu2YXkeNq+EoJyKTIegdSGzn1TY6pBdMkRA7QDH
JEKQJ93V3cJZwEFVTMAcLYX9oDEev7lzaiUX26AduOACBA4NesVPi2bJ0CzzDRBYnmN1RTAtLSo1
VTSC11txX4cUTcVeYf4e6UMVhHN9MYjZv4XI1+1oXtqRtJQH+nzEoDgVPqpt7zoKSNDwEl69scxI
D31WUg3myGAa0qX9xb7hWcvso2fOwASPS9lBreePcLt9lxCv79nYAEC3TMg4ereEI67LpIVOL37z
2S65yGoKIbousdB2qePzI1YOEddNVu1n8A/P31EmGvBvkAFbHpj+G6DpM6U9ROPggF6SsxZkKOWE
Tre8aKa28OqZxTTQbHpWtkE8uoJpNUeB9zIYBFS5+MyJ2XWRW/2jE7k0wh6A41PJGGQODHtgw84/
CWFyPbDYRY3IIbLF02CGM6cRHITkZoBNNLFmdinGnFMtWg6iBOAv9LeRz8Qo3onA1dEAVfbinx/c
+pcSzauzYWGoe79joY/yUYkpjryjsP+Ro3ZsljRRE97/Yt/VTla3VtmJmthVVzeq8+kxv4SEQIYh
rQacitohM1+RMyRbQHxfIVR50HhE1gxYdLAZ8Q6DGPQiDebZ0o7PDaSavXjxWS3bJsPgXT8IatDg
wkK+N7ktejuMvVvIAgQcxqA6SNrYa8E0l8ZLIXDuUHnM9BQjJLJVa6p5A/dpPC0EghJtaDA9qed2
BOgpuXPJ/aZUfyVVbqxPTnbIWkIIrYWGq0hidkotSkFu+VhS9E47219OO7CZnvSLx4UyakuTTTk8
FSsjBUi4511vJCb44Es42wzqsh9GidDqJ5f60ZHvhQxPe/amXyOFQg9LytQ6I8ihYqqAl6KA7tOa
pT/3a093TXe4X1c878dnu9KmXnRwDrkZ5nTdBS1foMAB65NLFAJ5hy5JltFgpdB0towBFwVR/1dn
TZn5ekVa5aSd6oFBl6zUzNfOLUHAnWsi2adwJ28ZlYq8u6MBMoYhj82OcV2T4939TBLWK85C8CfG
gN1tCLqVuuwcsX0XcNdFcsxfzgfYuoag2aHLTd4cD6KTzwdE4oBujdTX1wktLX2zfYzOSpJR6WKX
gHOK4mq4kz5JPcuIR4GOHyqaZFtKCBRsM/CaS9NRvkYlV89bVeoJw7+to8Y38symxoMTjS/pk9dm
eFrgIkgpQuoOeXFVADs9tweOe9wv4RAZUqB7x4e7b6xOYL0WT6/t9TEkO8ogaDPuIFTz1mhZBQZQ
053sSzaTXsRxYIi8/m3N8wA7qnlFLYEl9hMkozlv0dIi8wQOh/VQfmEc8OlbGDp9NagSsVytAkc4
tI+8ouBIXXjkrpKJBdauYXmA0KHgNE4545u0qFN+YxXtzY5NFklsr6uOJ2WVF7X6Kp96eVOZI7CK
VKU8r8l2/w78TLKp2sZyeKikq/ivl5xtjADjRgEGO5NHjCg/f2S1Xhcu+8rPYW+/SGV7BpTW738C
7cIwsMf7IL6cD0c7ZeXCKR00EX7W1Weo+M76rpVNAd9YSQJxUCrPhK07JihxGrZk9RxZWe5gVWxH
iz7qydfpD1EOXffOAwECwZ2wzF9j5V3Wtj2mUMtQYrOdS22v6MJ2utQwahkT4fHky9wFVTzmImrf
xf7zXyEAmpP58fkhua9uoFXYyRe1uaNB+GJdWsppIltcUppOlO9R9+5BjtMlQJVhXygGPzvBEFef
XUsBdK3enVULI/7vs2ODr+N1CXYDn91GvJi5azzbV3ZEZ9ErU0STTOwOiO+Ngbh3Fisz7GUZm99J
BORy/dKVWAs7MN3CXDIC2o35wQxvlTuG83ZwIsNZIWpZ9Rsv4UTn8viCKRP3REmRa7ayJnEzqj73
aj+ONXY7jsipTkKb+fGoas7yXnz4UFjOVS1DaJAot7gJ+pdbB2MhJfFyWB4twQgkEr04wenhhfzD
XvzJHKenzrKkUxRt7PRnBDEamcycE6oLyzqZOMGZocFui5IeFh5F6+JLYG7MAZTsmV4DxLx2Lir8
qAB+Q2jCR1Dnj+P4BbiOo1amSA1NfErFc1pp5QDu2o4tVe3pqGtHjVein5L1QZGqJK4ocrh/jsR6
JiMdw76X04bEsw/N86GDCiGNdzluXLCmWvGHMhcZo65w4XXbE+1hDutKZkkLay+T9UtVf+r/jVX5
fqN0yszp0VN5KT3EcO4KoujmAK024/swU1MygM/TZm5eOIrkSbF3JC9bn2LRSYQZU6ni39pcNRLC
gVIqBF25SUn25/9SYjYq+WrPnk10Cyt6lqW2aT/NraYjlxcFcMB9S+LPS/NxYpuqHbaO8r5WdKz3
4siqJ8WzsYm1KFb5gZOP0Ofiy/ziwEZ7dfN000/Xesw/k5CeIh9F2Xv3E+kCtDYiJZYLRUThsY7P
hA9Dq+Put3RFzp0muSNoLo9WlZ95YV1SWsw7AkyDR9nVQFR6bMBRFFtsWBu/ty32apJ784UUAzHH
u+G5nX8x3eOkHlE8OWpda1oFrfZOBK8FVj+LrsK+Vvc/rXJTxmGRM4mpNZeMHFp51Aoi0dutFuok
ath5NpFbRuamTfNgw3j9eYKYFI6Uq8v0cQBKkRyEN+bcrtfUOsPYNtc6YnlZs9qnx1fhFYKKhOMf
SFRi78e1R6qlc7f8VgyyN5UA+HkS2yV8IQ2iVcZ9X+MKtJOVRSOjGtABSwbrsHikS9ePa8+lyCrl
OdkHUknQRZaiB9B3YVKRUwOQ0NLzapt/ExwXVk+xGmW0iPenbJBwIj5s5E5Oz159Rb/vEmgrPDjD
m7TvJbgbz6/8nTWsgikuyVrZSbRAFKMyM9Y14AdhcPCJHIZEvtt5IlUoRAn+JXHV5Y9LdRt57sDr
HsL/y0l2bAazucIz0pcQf906X56A1gGSqUNrtNmUjVkEpsiwOD9N0e0R1R7uL536UoVQt02jDP5U
pn1VgZYPCMzlUvPUGtl+dKWoEJ4GBaIb994fyvvct6rrTz/GlLkZNTwMYyuyV+heunrvGbE0ksyi
5QAvMnc5yOOB+1UFMwI3PSCfXidTp1Emzk9r5C9RuVFXlR+UtGKUegxNHKfGsG1q2Czqaear+SCU
Yczwt4Pe/ZufzoUamdvUFjWLQ5nm6wZ3gOS3Ap+jb3XK5U0OsAeOjbLSKTq1LOYd/V+yjpBuPaBN
+voviyCBuGuqE3hmFfISAZ4vXMPu8AXbzb+RJ2/o/GB1KWGPHQ73POmfg2Eo1z3Rq89dWcUbHDha
zfEGc8h/iG/9jDhV6zoTXqNvdEg6XhukNoKdQ+j/Fa6SL8g14zJRX+aUU0rpuKNssadCLKnFDUyR
fT49Wroa28LnHnMNgpRZmvFQNDMJaeIqWdGczYzu31fT+399/796+/E/eaavVu2IJnovTwqcVkuo
xDCnbeeruQRIrb4MaTfuWDTHJ20N34WmD5CBjupNTvgt5qIygxuzgEDtaF/SJvV4pwQKma5rSzlE
r1s+TT+t0qQJSQdDNI2C44NHIqSzoHKLf9CTMfsNbdKBlCKPJhB+VVl50msel24j5SxkOTo7u03c
I3to/AKmm8W2rwH5kQ+i8yeTkg+4lcqWp8r4Ah+ibFa/+v5hvAMrEoLY8gctGXHaEwKIaUU9jipo
jmFkjIzF3lQ/8KGS2Z5rw78oTDCQZda7u3DKFVMld24gWKc5jFibxiCFFIDMIdqGYauLFjLelTDD
lK/YLI6byiY1L7HlODo9eMY/UH9BzrsJS/jNKL0swI7GulqgF3844vySE76+O5TjyXl219l+g3nR
TZ6hxg0gmvAEz/KCDqHk1nNWoUlxnjvx2qiobI8cXrVtYj0dx0rrYu9p4Ug1P4LKLOb0N9lPFzU2
fjhA1S4tTi7JKBqS/Fn+TQgQxMyXPUsxdlm7j5E5ulg46b5Vu2jnamrszL3Rt2jqg6vu9ZDpaTy7
6VRTwJQLcRWMAyrp2MKq34Zz5ix8y8On0/lksyAGiWt6WN4NH2srbrqIUdTOjKbdM1wFkvPP2azk
wrlQwk9fhGcZJ1DkaVo//T89iUDCYowNkiKvMBiA30mmdEZ8wWVF8u69kQXIQOB93w1Y3WtTSfpK
Hjmblan9uFGGCdyVpigHSLHcgHXY7J8SJvckcCWBKaXmzUzRfqI3Ss2fwWEU+sjmzGd11HfeDTys
3svPdgt8QaxacmDvsk2FavfA4Kwy768M1ocz8TrsQg+hv0VCMsXeVfutiFZVQiYmtvj2UCnxZ0Wn
49h4W8RjvW/kMvNjUKfQsmuPicmEhlqA+8mnonpd+TpCYgYar2KfqrstSjwCT6/xsup94of7wJXJ
00ZNiYxy0VuDdZvHUWokpXfK5NRuRLJgxxgt5BvvmJBEl3HKs8HnWp7iquoQuj4mDAOpTFzYFr6T
z8LmdUSSA7h56N/MMSqNCX7Ahe5sZc9aWRjE7RLuJemMEIAoE9z5SWSFwQXbu5y29+QYEMykfa8l
mY1LTQGQ2LAVQVgIbWBZLGjcobQ6orh087Glp1HFAh1GrE9B8LCXyRtYbCnV5sMmeJQ4OhqmzyNe
ce75klB0lVDJx90WqS09XodXA65QqYo8bmp2IevINAnAJTywTYEfW8sy+iTaN8OktN4JE0ir/eTF
uEPScevYa8pWAV74QMGDlx1mg/WyAaksdRXs2dpS4L2qm2PXzOgG6X3iN96UuM1ReWws1BoYonRu
V18LcjeII4SokjcaYbZBExv60N3oW5NKkJkM1LNsTLNTpgb0x8SsotFNsQ2L8zwMINLZYumzJSqY
uCJzBq/FPQxvwLsuhueJ3a76otiiSPl2f93fVmrWqmlHZQ8w5LZ4QyfHcMshKuOHuCSbEQGokYIn
f+kKQtoM0+fK+8/Nl4ecyUU3dwiFqq3CjDNy/mrmGb6A9WJ1Jp21/NmWyzgPEFtdmSXu28DFHvPT
f4OKDMDpgZmLaBW2gtM/gc3RNclFCq4s07mAGPO6pAbw94ljpltGqMfhX6w48u1++m1Y6ejcZsNm
SCJYsjYzKgxGgETplxsxU9rux2wB8fqgDznKoTkcBSk+21vu5j0ETjuqYAp2tjMPsKlNqrGLSh7y
CnIVB69Q3XLfMWY9D/xzus/O7AnAEIk4yHWXGIilCcb0eeYzrKMB5gj8vOrEd6d0lv28/yHxEdzT
X/uwdc021EFKTx+AXA35JCYWzFgesgQfjB/cVEqVzdppXxFOf4MtwKL6AnwQ3pLzobdQx1FmCsE/
Fe6JV0tqglje/T0Bzr7TyxcpRjDYFDB048oKqshtQoNxD09BqrcNJLtygm+Oi8h18Z+C+HlMcMDI
cMjRzR+Syi6NeMu2JNBj05lH9yNgzNBzPCbGxXb1hqOHIJgpscSPkoi1muQ5UHC208aTRhb8DDPF
XqintiXDrDrCnXrobdKFhGgfx8lS7BzCqVxxWLqYqJr3YZCOHsLi42G1saMiZqXDHWsRfcQwHDsP
75YZA/nCtu4FhnLQvSEtObSQU4rLoIart8lpKHROXBkJ+mR3XUbVwGYcIKNsqUJonfeKLok8ZESh
fvS2JRV+LkxFEc6PKIysA7WLQ7mq3nCMwFYI1DtJxfRnicotfw13NyaR8p7bdlnENVSQdqGvpLy/
lEOqXe7NjuHnhGO1SlWkjvWt0EeHilwfQehXEV/d7/2PTWHRUhTzBsLPq8Qw5XQwrJGCUkNqsGo0
n9GW/1bcXrlSio+kf3T41KlXRTrZ+E9AaIltkW8q3nJWnyivAk91wyMHOi5dcaVvnO0K0+myuEZ4
w2BKmZYrl835hsjP3s8bCfPaTE58qE7uxWv3Sa5ipiQDLaKOyKEl59waEyp6cpeRdGzG49Xg7QNl
VuA6p806Qf7kUw2/SexjCiQGmicOSpQAVhjzPGoFGeBV7qyZSh+XtmkpvlzgazXKR1ZLZgm+cqe0
etQoR6nVYwqJ+5IhuUsSgn1bKyR/hcmobs7Fe0ZgKo+yOw+vQFiiSEb6b7hsgvTehY5Mz/6ppz6I
4Ab8RuVrkGAoHiz9dhNe0c8E9Bc0QrQ/HkFFu58dD4OrQizCzguHZ1ztcxzLFXDcQM772XnI+b31
tv5VUHwB6puPL3q7fenRR4FF6Hq04mPR0YpMPSSMtsSzFsVI9XiBzVMEJYw/iXF0CdJNLBwjHX6A
2YO5NqF34XiRRFliSSZzPutwdjo9XHYYfL7j5DnJHPv2rITerxo+TzxiMjyR8ckgam7022dLJKBK
bCfFxXVNwgx2+59MHsYIovod2YavduyZ6p1Aov1tYOFaWppsEPArlwlkUBMbCyU/vAmLmpDT0qhS
XAXdiR2ybGvQzMi5D3va5J2f4hg19Tit1VzEtG1woFuRzkWny6QFVv1FIlSPj6xgmAIxIx1OMvU9
ukTqAVQObrclcqHfIvZ73iVGxgxpt+BGwywTZcZltygzgCnvO83n+EoXdp7PR7Cfb5Bu07M1Ujdl
D/CfMuurkxC1xqSLEQlF+EAghXHfi7KxLDEgBEKsKjQB0OjYjkHdkDIGyIUkLkgQdKks0qmUSDmf
0X/veSEagX+RcB87b2qIkoIeLOkFUDbm8jVi/+t00vFJec4ph2cO9ct7zNYHxVlEuyMkB8Hxr1MO
zyb2mEx4hJxZoSOrrh7bAPoy1Oz21ix1GrdSyjzxFdbHIKIZUjP9iZwlN2UYevfugpzN/FmeuJ58
DSbEFcOEJ1dLTOHe89yxV7g6h1WVVrPRiG5jR2OLo5bh9coI5Vy08wPshoT3BhRvQv3dIfsmkQeU
8DB0Dq3u6RGDBF8CD9RSnzy3oORRzHmH4SWMdUQNCMtzD+ljNjUEmQ/0lV+5Qt6MjDShUcahQIk+
gj+XbzXPdq/lj4MQV5gxzDmX23KyDK6jO26vRjn0jUi+tORDR/0+NUncSEjlHGB6pee0vgv/BLUl
HFdWNGvzmzkwSaaRBqqrVbQvUjhWOG+C9ntsvSfevxlBvv1e1opQt7001UK/0Ne0TR8l8n+mX68h
q2YAWCGw3lwDpjWwn33DxDWbEujpIvP1cG92Mf/fR0C+/G2k5ON3jMW1Dy+SOOJBDB33rV5l+XT5
3OIauvdBGIycSaObP5ilUrva16mkaZeBYivO0R7Po0zM08wiYObGBmre8aIZnNlm9AxuZ345NoS+
akUEjAbmVoBHvDroNgE3qepYib8rRwxQtxGUXo2nAKwEehnTCvMPq5Qg7zfYq1qufHeavRRmo7dw
QEKkhgJO+1kDTpfdSCMFnfhztN2OZFYYUO9DRt4WReVL2f5aW5r6nIkGOAAz9bYB3RjxWHGwswOe
Wab01eZBCeS8+O2SH07lK+Gs4hAF+hn69dNugCCWxBGiFzOf4SiHiUenBjlcrutrPU7gokKJGFFg
WnV4Sqe00QvD8eEJaYRKNZeXY7Wg2DfREidR+sfsf7nSpc8P5Nwu6VYKCLLJ/W5ai6/auMpCfyAX
npYsEWqRwuBhZqFRUSNu/WfuNqqP2UG2hmXA76/HxLzRsymOwDOe5f5qLBBIBO9t+72aP9qx/2Dj
SXXB/UR82eeAxl2BqlSjaIEZB2foy7RU4clYjEquyXPammAvkQWuKrqr62q7+GBCEatHfGsDlwF6
lG/GNAnjm6NTo/bgP3jxKj5CJrja0IknE1KObgvOM6OHG9c8KvQeGXKNH/JwKeUTtfV62h6tJt4b
7+yY1q1lhgbgBngaQINhPwNXgeJWL8Va2uBsmxIYKDCzqiaOaCAH7QeW0YRP2KT15h2zC9VHVFIV
JWWap0bjEfLRqFAdt7k0lND3W2/xR/M10Kzyb+ZqcecF7kx4enbKSnTBppE09Tg+0CxiMjVHL7EA
/4goo3e+3cgd04pChPN69uCuSkkuYxPQM/L4ATQrfDeR3TwNiw/dbSAUaY64vfxn/VSYF1YS0htx
mvNIPH1cb5ltYryp332Ipp4Q+vP53lBI7jqF8u+TiCwPKt9qmGoO08CYjpkMOtlOWRBtq2erfkWG
E62C0brnZw8OaEFnKaDolW/zzeM5ntKghr8Mme4MZfZE12cUQhmAd5UlBTp5oQzkJhwXAb9PApCs
lCSvp7M/0oV1CyRO/yiePx567jDOJTF3VG6BiN6nTKEi+FqVO89UcN2+z9g0SJMCu5n39a4c6WTN
FcappIn4wAW49Gzy96PHC7BBz5gI03e0mNsNXijj0AOyej2LypWTSkT9u1rQOBoS/Vvy7cqAXOyv
/q5gMIFNaBf4aaQmIr3Z+s9Lvq/viQdJnq0n0EFVSDjzkJeimZ1ZJQgVkbIY0B16fN+SwIh9auQC
+8key4V7CZXQcogGdD7K5jPy62yn4SjyOSwdFAT6zE3ZxkyXkJhEaGTktXZmyAZHaUwXcBFCS+dx
GscDyxF8ZUQGg9zOHE6odS1MYJMPA8oR1fyI0Khqcw/yUhTkbH6wmdN+jzZhvjaydurlHR2y+3M2
1aX8esTBBYwE0Y0E9oZEt8+Cv0XcGOySu0JtfkzDk9kUs011bWOZdzZG6WSAw4mfrtIBOOXiIYIB
U7SixHjWhaZUgsi1X2MuIcadMDmXzz5ljAE6a/g4OnvzOShPF5qbI4AarpS1OodElRMfyrqK1B+D
Yz3lMHPlIqlrW4dgRSXMOOvXQBNfO2nO893umh9zHS6gKKbwwsh8j3w5fLNODRECNFHCd7HrbKbR
1sh49/dDCVWbTf7hFa9Ig0dol3R3cMiWweWCNQi/nUNLbthc3YATeGt20wz2mSj4GfK2r3RCVqPw
vwyxK91yMWqZV4W3J9hAFFZGIgAFxBTp1/qQxY4+IOv2DeV+HczhZsKMxggQp0Nedzl7SXoUo6Ym
tJ8nHeW5PHcgCfxyvDQ1H0ZsoL58QVxdheCWOq2q91t0KEI6gs3kRY5+0VVPAtUoQFs1heviVQ7E
/t6wAUBtTwyBWNBw5nfWu/aA943wkhZu8k1YVliwWUhWNQ0MU+u1laSy7rxFTP8J9l9iEZaDiATn
jSjrG9Ryi36OBsTwWTL6JZgrOR2BZMrg2nIVxWcwwXyNeowBV3mVWmUGS8qoy6k0GXzI+x48PKL/
IX3m8CV7HIa+/sCHXxATM2pqx4E/7EdNE/v5UEMp8ab4zgPB5b9rDLLoKDHctHlp66pbmzsGv2S6
EWElNna5fRC2P9dR6C4sW93eQ4tT6VViv44YcuAU2C/lEIehxvqWAV9IQ49Piz/taQJd/4mQq95b
QyL38sBdRT5bTMoO2PWe9F9xmIkJ7Vj5/vJhaYUmiuq6wXfGsAVb8BLEKn8Mxe97B72S54UCZGYk
se2tORHZo5JZRWChLV35oQwb5lhg0Ib9c909kkIumQzGjmXHOhB5I3Xe6aRrm9TO2xXCXey2nBP+
s6NdzQ/KrxnAdISuR1/HkFqtC70xcUMo0o9AXIw+heHhxUV28BGK7axaXPXQwgvatHslxTH4eJJf
50IgEVelG3n81sqJdxAUh3TKeDOK1deL+9ErV+yK+PkkahbSoc8LUv0XyEAVTF/39UYRbk9RCzCS
R3dmJLiypX3+dK0sDPpsdKxYu8Xn6gF9wnA4yUiGETs606lAghhpKbffDcLGUy76dcflD9DRo0c8
6AMxAl07+46nG6My6ZplHMrd2HgmTC7NJIs6RxszV6klVYu7oeayqOgZkZBdiSc6B1s7G3Y4uQ0a
0oE4OuZZiLUXPJXfdvNUNIHT+P32PXnHOquv6g1KP9Crce85ShDyZ3z0/2MXvwr6FYLiturqMN3J
2OXm56NTPLc2/eiFtH2GL/obF6/MRMajclIqUzKqGskIQFrL44ke3aP+7lZeT9IVO0nGvgQuH1ox
eoHkguB05ZWqJZtAgXE0yveKff4XPGQDnfiCNdBFQazqqDgapbqJ1tULIQUnhgo56lg2C+Z10O/d
72hOXWVPtkdoGM9dHr4R9+mr9NDZLHcHVkQabi2TzzJKkcDAduiF0syw2y9GhEmx/X7nLzan2DVA
EBIW9jqMrLZ+vr7IPPgD8bbZjh2VCSCf4IcKo08IbjvGkfpYUrVO0MTKAIUgNTsgufALMDIoR61V
M/7zhU373FskNBc9xe60ITb6fUVN+ZpcLEmwWzG73bN9w7Xq/KLvG1o8AnAHV2/vI4BT8enFSFY5
io34go61UrmT6M64zDfuhgl8hsYmaW6Ux3cMC+BljWsBoiI3Gn1UKsdlqd03mTuxrhurvw5x9pBZ
1ryax+yszIu/1EaogoptemSeC3vrc6+ZH9uxSz4LAlHFUR5iwyqmvlcdjSOcZn6XvB7IlnKGqYQn
g4YyWyYYKQVGO/+QVpgABobp1TLDldJIAXhurBtG7h0Lo43KRtJAHdPcdEzm3Rz8dCO0JbwFZsqd
REbSCidkiwJ0xC6JxvMVgskIoqW0f12Xnoj6gDzNX6M1xFe/Q57/GsvCbipZBQKV1F3aptiIDVPm
5lhc7dlQUUzQukoZKZso2THXzwSzT3Y7b81RuTZGmmwX/KB/CHtPSPol9iT9T1fQ+/NeOE0dIInv
UlTve7LAVPIn9HsoR9pYamo5rq2jIcOWUWeuhLVQp6bNKq5L0rxlbfuH43EXIb1aIPtuzviMNx6L
q1Q7IsKlctuEw9XYkjkUHU6OpOzQOFc8LvHKNLZMRRmiAS341da9SClwbZM2OZu5cTqRVO8c9NoM
+iO+cQBSjIVsTJ4A6eJ1cC5boTSS/ql8OGC5q5KPIWP3CeECwDmwMGK3o7mZeDZwu3udaQ5wYl7p
dpMtbrtvTrCbq5TvsqWkYQDj5+VlAyxPxVkoJd2osvghvE/puEnNWAyxzRutksSqQ/+4hPRMu36v
I+DK86peRqqjd2dgEKjufAmUqW8RDzEN82+O5uSLu95d6Y5TijHp/+x4nHvi4noO1zP9Ioimar6k
XTEyx7sTbRKfXNabtw3U8hyBLb7dhwfKQrQzN3gAc1uGpgNjYYoWFIQUBvfpdq/SbuQ9aqOQjJ6v
j1TYeF69e9VMoh1LBku4PFU2zBICLN/TZnHFL2XmTlTYj3w6xdTSdUF8U9EYdFyrvC0r2rnk1HhK
kH9wbBfxY/kRRleoAC/OgwUSpj4/v8BxSq2kV9Xu9qSHWhD68E7xUAQUJ7rGvUq5LLXv0Lr3ML8X
ZzRocyzeL/pcHZ+V6vyr4WU4gLOy+i93kY8XiWAjizA3tYY0cfG6NDd1HsyV/DFHAcVGeG0+QTUk
myjGPKoo27YQmNWD+/RNwwi3ycJLJInK4BV+a+FOXPqOJJmfE5BAD/uZOufUjYzwLh1gzOYAP+9R
W9wtZI6/DP+oFywk5DRP5QZ6naYAFUHm9d5OcTLtES1mWAxIgJvN1T2vLmiTYhjkEqPuJdWy6HwD
MWeBxTuEskeG9+j5OVBDOUBPPt3CdbAcChKLkV2313Bl5axo8wn0rPCYgR/RUin6TaDE4hzSmEDm
I1M9s3FGujdAOuUZprLIbIW+L7AER8gF3s8DtCYjaUMV1il0tNp7rD+cIMpMERscejNKzHpVK0at
eNl/imDZQAAMTACmdrCqPalSSa16xDP9ASePobXkvkXcMCKGQw/CgHTULN2Ij3WH+0R97Euq4w5j
BJBpiT9irZFR0sogEKhM1FC/lhvrWz+Ag10Max0WR77yN9ibKitPWpY5rN6NM3tI/ny0uh+bByhx
zJqLtzuuTPe9+WxPwVsmoRlMnIMbQBJIbuFPc35qswS0sd6WF1YOmWDoaSXyKfc1AAn/ivZmPm3m
tCofaRHwtP6r3PGKoK1ozcwfqQ/bROVx4rpwkDrIk5+VDH2COMvzEO/l9pNaXNTJOPbSyALR71g7
rYKfyJ7FvY80ZhLrw9Pc/WYtt6Fv/ZfUpxspf80W/ltD6fOS+sMIqJi0ceFoCHEbcRoWHj31dIir
sQIei6US5lXrCLc2zruvlQiAZ30E7E6EdRv9x8j0A9vD7M7T6nQ/9sIni2jH3JQ4vvwVhmnigWWg
lQWtyxY0WbNWv1CUmA6B8PUx5MLw7EG9uREmKcX1ASgBd/AgmFjqhp2q44iBFrJ+csWwpZm2//eA
Ij7isXMZXBMj/1eoTTj0r+AHOkMrbHhSabhKIgNWd6KAY904xzYiaurzgmNxan+KtXpERnJWQWiX
A9TpZX/oeRpftNo9KqtngG95BKlpqo4iFnCWOVUxILdVdFgJEjVt/eohkEfg8flqLWz9UVB3HKmR
qQxnS8SHqYW9hgVSrFSqZZlO9YPIrRBSQS4HBNdHO2FEYD86fLAPxvwbQ9k6vCqe+pB0oqfpAN9B
3N0IDwjp+kZPvAFil/mOm/2FKibZJo7uP/fYuJWYCkj6Rzn36fL+G30K+d0ZeDR7oLw4Xf7WITsm
zHNscc2jVIfV8U0L9gYz5umgdUUk18WtFaXHaQ5E2BYzS+BzuC4e8MrrFmdTe6rPqEIs5W6wDmX2
LcZBTsyt3L+FEsNDCkTMzE2LrsWuiDfjzQjVad7DNHmvoK6rN9xYH7KuD5gkmXR4d/oi+G1FiOfR
FV8epzYC2hAwzebgz8Ky15QS6TVQHak0dWInPYusEiENVvlFPqkc4Fbc6FwH3bIFpaQiDdE3OVY9
TVarjeoVf7Ph/9dAIsUdkJLAS2MiuX+KQHZheOwY6Ui2NI6nYl1CR5M6hEcwb+FOmwrFMD3ZOlIi
hwSh/QzcbVmYx9H4cGnbdMIa4/9gWgJ6IauH10T12G+SLRWbvM3D2ETKDPkTcAg/5oj9RfYzW2cr
oI8nTgCkNCbBsqkAPpnzdgAQF0ez80UGi+VrhrEtvYwScbO6xqovHJ/CjjBt0E/WkFICVvv662Vo
S6uUfhrKCPalcIm8FWSgE38e+x8WFzl13nIlHOuR+R3tW2b5iAIgDjwX3z6BjPClYGO1vEaWGIig
CN++R9GMkut4kwJJ7UKlr3O+tolYHBRvfp6tn+BxYZhyhMbfgrWZxWS/5YkzYE792fuZRDYUdPqp
gLzegd9IceidYwriCvWAeWf5qKm/Fki1lkhOLBH9Cllfn1F8rLt7xE//KvrdZwGh5P1Oy7GRMDFU
rXBoPq1ypbpys6Yp/WgegjTMCcRc2h84qlAub3eAeqID73o9q+1+Ttg6fJu/hTGGHjZJYcRjLFGe
EteBh9eIB/Bqb3ZZtbxIoOAAQFGxSE/1lFSM+OR9001DNjTygMlrsMcpxZeWiahhl5YP35hFNDpH
6tHsFxdL8PCziPsxZUYnLVy6PfPNx4WqPD7f4otcnAPbb2qIWSe4r3gvX9xWhVJhEHFSb6IQAwiC
hnkLULlsv5qtXnOtQCUoNH9I9FAQTfsFsENHy285H4JSM/vxbqLZ9XAHx3qbEjDys/P+VAO6yU+/
TX8LnR3ywjBbCL4lKMHO6SbktOZlSzsX8tySoBjZpov8m8fpBuHBJ9nBAyQwzwFEYCtWnbA2hHdF
PZ4wNUxfVIQo7bMoZ6hHsplSQP3BhhUhznNkoMzBS9eggz8TpuBPgSCgCkho3hW6XuML53dNQWZ8
m+lW/cL3ZxdC33nDnEu4QTu2kZDHqh2qUw4X5e0Tmlkz9ocRrXbqLPq2bBDede3BdnO2G7ne9w37
9o8/tMD+uhaf97Pi2qP8FNudn+Mk6DnLOAnReNk6T7FvLC80B2y+GeQ/6odkGevzfSGOEwV0RLqd
yhMHSZp4ndkqlKRPM+UZf6xwSHIAMJfczt18NJRnqkKZlNobfsc6uSGBlSKFO4zWOXrVMKSvJClH
x4O+5VpF0njpmFTozEmYE90Kbd5+oM8MmrvnoopEuF3HuvdTkz007X4TMIbG2IdCTIlPhatI67dm
9FR8ztYfnBr7qt5p9YMCToa3UigFkU0PGmGHmpfo4Df+H1sb/7j9nPShknrJOcVDNNErLVKzMNX1
w5BeW36Gmj+EzJa8wF2IRJspHA/buTVRRdIsvnI/l18N7ML0hqv+2vxvMMz9Sq+UQWskOvODh/b5
yeWEwzkfLHokHfevtIlzCOBL/NflGZDZM1f5DZWFIIHIsPRK5tt+6DjRlMb88tSahLdPdLkHp32Y
MEfy0ovDagxwjpD0rczBIgHbWenrLqkAAmxoo4GjaHp4wUFt82ABBHvx2rQwmiz1zUMHzHkdVbs0
0fa6ovJH0NF41YP1RkGq7EhTnfjxaVgSyysr94rFDTr7hJHFoYQWNSf9UAaCR1Tb0i8mzq637JLj
/yfGpooVXkKD8eou02pXhPfh7EaO9P2vhyVt5n0rDwKVWP68SvLwyAkpaTPvOzqJgSQk9tpeRRyS
j1Wf/Yeud7amjLX9A/3zKGGjy6AoCM3e6HHADPrrSOXZyic8DR8oJyfWn6nEEhIJuTcL6J8T8GGR
4smq/Rq4JLQxSNlynDquXQyPYqVcUfOeFrgzLpvfyT5M43qZZLSBO1e6ukua0dn+8FXr5tKfv0bn
qLRNzVM/PTx1Io2s2cI70cUkd/ZbS4MjyajTJwIZAdKMaCmAto092y08pKV3yrROXb2iAyasMw3V
9ijQFSAd1fLw3vzaC8jR5/XG6KnY0UShHAcgLIG6Xn1IBnyvEo4yQ0jAV3pCWlO3zh/dXBIAzI4T
u26pzHTSm4GBC/Y4RVjqFK1Xu+rAUX6FCJNU9k99lG98TfiSxQh22Vtro83tq/qwtFt3DHWkaIUP
4o9Okl7lqrtN7rT5yOm0Pq180u5RM6VuK358uaZTL5yrZoVHLao+ncKkzpCfYo0Oo1r1+ZdClmf5
Szx5blF0DFP2Z91vBMom9HMz9iE4Q4ioKxUek4l8ydcPy9uMOP8DTeO5xdDgDk99NSEaTqwHiutW
/QVek4BlVANRPisPrm5w9/mb4Ajr+1nNtteI7EPEKm8+lGwXENV3IE/VFK6b9C7u+gMl3OK7NhJh
l6CXoC/OQa7K1TeYDZSABlUwMUjCAL4i6XiSy/eb7zENRvC9l2OLJJ5vB3tDIv4JxOBSpQz6c4iO
oJqh1MAfq6Z3S9U1593KdIA0c+ntq84/XHD3h4tIhsjt3bN/STGlFjlquGnLDVjh9SBzl2/eCb6G
gXVnxY9UcZuHh9LzFCnIIYWzRRnnNBaLEOvY16q6GW8gsmK1LMDPuXV60CwW/HSeFJbM9xn5ff67
nXkcCs7soUNyfUWadiFJ6T2PhHSiuQa50vC/9aZRcLayhDqsPbzwLJcMItd05zcRkyThRzFCsCfQ
0RAl6bhiY/Ux7ocKo2Qfmkak/yewx95asug1tvFT9PhnaVAMFedkWaBmzDM67dB2qxTNQ2Pbzyoy
efz0dv10u2KoMITZuZHqFKzxr0p9teAUGEg9gGHAE1LGebHLYxH6oFkK6zYLxzDDq4eFg+poA0VA
Wrflg6nstVy+xrYaRYTq64VsmryEaZPOgbguV7TlFdMOPLiOYSlQC3Px5P1PBl+N4+dLVOo/tY28
s4eKD2V3alA5Vu0/TwUm8FvBWzPqCPy3e8vPOayrh02zw0CnSw9CHB7jClFYX57xYA+Tv8gYVgwZ
/+DS5CherCS8uBs161tKZu8EBNzLAL2d8AHZApGRvBNnwROmhopznMhcndiSXSJXAEEliHileSu4
C3ta6LsCZ3rY+vH5Rh9Et/MKjGXM8CEc2RlAEs+4+RAcgNLdjOnD4wELWQV6cBBl2yWTz4p28yV9
BtkN/O69m0fDj+hPjLpBG/c6cCJLVTeOe3BbsD1/rIrx8S2c1Pd85sj8lQZy5RYFACQC1DfH52dt
jpeciujX9Unub9nLpj9nq2dAoO3aXrE0VIksQWXK/NVy8vfPP96PP3h2bHapGO7LwuQCJL1akLjG
tQ6Wi5MH057/YCldEaboAfZSG8kQGQzdnGA4Ech1Yuf826oQ1pykaNShfdartcrXaVyJNx0mlV3l
iOI8NnodWLR/2tJKQ74flS1yuGnE4TPuNvCA5jmrfkAYf4Fb22ECMin3rMQGtTgy2a4imUf5k7Kx
5K8v79wYkBUTHV6/nOPpPqc7xUAHf64giLq0alFTBcJmSeK6cwuLxPcaYbzG/pgk0IaYBLpOFYpA
JQIGa8oFaiDcawtiisVIgylNCfNin3n/sn1Yz4dnVqwcc9R1qPJIcoqfwuot34aXpk0YA6ZLnIHu
TnXSj1Lilcy1t33zIn2cRoqdng/RZYb/XHMrg3ESQHCKdK0BXkv6hk/M5RMsGpVEtLrIik5I0F6H
xO+RhpFGHuIzqVIwnBIgsV+pi3v2MDf8G7jV+CCnfmfxaeqqzaQ8yZt5/vzx++XAJpUWrDEOY1Gg
2UMDH1IVNRZp11fQftZKLV8+3U2OK2fLfeDfvN3HANU4F1BFKCmU7WjH1zwuG3JSl28KHTghgeJI
TWNGDkAp0oSTT/4ODRfidvMDoWNqeM7p2vzlz7xJWs2en8SEDWDkew+EAIVPSQsWgQMx8f7Tmk3p
2TFFH8vhSXevHCdHr+PzQM+T5BLoGLNTMp1de7V6TjK5ydusjJ7wbjhJ/sH/6CFIHgKMMhE+UJai
n53KJMJlobGEPv+SiwbJMLXwueQi4lrdTFKW/K8JFcbKq1BqVmC68IUZUJIwEG7XJg2xzwYr1ULO
agdNykRchcxoOqoQ9COKZqRHY0MNmZ15BhYVQzZcNaG7UAXPC1sQRvH5a8E9URxXNKqbAByqFYf3
c/teFGVXAdG8BWYVdio1+JDUDb6SzwBX3x77QY6N+TOCJO1teUSNf8zCznf/YpcD93qD5Yvmakxq
8uyTO1xdfIoW9QBS13aypslYHX+jA00zgZoHUjjZsyDAR1hn0ATreMvNi1rEC3GiH6soTeQVXqXT
WcUyNS6qjVcwY34pAzgc/DRQTua97Ruaakd5UOac0D2TNQrQ8jEmXPgTz9kZF6+RZvlnvIGyWyGl
UqmQu0OfSJJxxBFjgDRodOAy38yH//pIIcGcc3jyxrBeHpcWJyTleZdHjqyJ1GSaYKlZeL0xsQ5U
FtL1clekvj9Gx3674vSNeANIeVZtytAAbjBfqm62f5qK5vq0/ZhDKSOqMR0HYGOPxKsG+5sZSJzZ
v91kPfuu3lm+Aa/7v12TIeiKAdn8wUddDOe9c2CvPFPhcF6kErIJsjAVbUL3gbHHGLkNb7uOFgKn
dqxxz2jAsuqTz1BB1WoiRuIEyx6z9k2pvQT51rrr524POq4fIR6iYxkAO0YbrFWi/VBO7lZQ4Pqt
blGC1+2TwfVrRpjKXAy37kaXic/9W9SI4iXvOJIGwvnkAT7OjmTnfywqdrFZylEcSRl4/b+LI53I
gq0t7T8bD69faE62PWqfK5c0eP5VNRHsZ2dvKrLu6+FcBA8slgKcWUu4Olf6LSe6ZxKrbjy2ZL18
1YtLDBBuEY9b13XPNClqj7orFX0SAXm98SycWQvMQCCEl0/q2pOJA9DMPl6AMarxjIywm1MjnBU8
u3SnJnCL3NYBfvsEFQq+/ox9tZMC2CKOa0XgekdsNPo6u1laO9ICOWirAgDJxJHnl2JtlYFk8yjg
y6Lle03KPLi0d5iUHy7Vg8Uvs/TbIdIkWhS30xE3NF+m9FU6GNbvikBF/429G6XbxqUBcjrGx97G
xPvkw2hH/NfXTw4Z1y7OyU2mqTBd0WcQRL8Svlj7J03Q6cPqYJE7mxlhKUr/BkooW3es4GggdyJd
Q+FyA/3N/n/3uFDgFEObYhXh83VECF3p6aePqr7MeR1EEOtwCSTckBi/N2Af+xuJOeWpkntsP/Cy
VKu9vl8vWFOeiDI/Tbemtuy+G0WAKeMWqWz1PrcnoHLpm2CkB3pPSfh5V1qX/Cx4g33UXe27MOJh
s29hip2qjLvEWIQNNqrAvGN0AZPN2x3YLUMl4RftQwoGyQvBTsgcHsPt6Q1MAlYZM+8w5Xj1hU1M
VcENnDP3Y424fHKwF/RqtGtJTG/zVs2jEaql9NoDcdR9oflEtWydCqhkkTEk6Uc+5gwVlGSG3p6d
OkeUrvbHf88WsXclv7fGZUxHk7ocaRUDOuxrGNi+9JWHSIM+B2KRssPJd8ukfSPWbJBuNQgREFqD
3/maD6zyCNhgihewVSjhL0O5UM0a0feBiznIRgvOzwFNVlAzj86bon/kYP1JeBmBd+FYvCnxLOsO
+GRaRkDHTnbXGPe6yI3yktwrxA9hA3h2+gsTj2QGKfR58c5/+c5w0QKXqWJIACgXuPVtF48I3LW+
dCjDOfbySDtV7LgsW2OLxYe3X77x+FV0fqlGsAEK0TZDWqz1xswBxyHi2yLpFnPdfD7QlIxHPl9e
KmziMCv1EoV0kT/cPmsV1pP8tUNUWI86fwR3/OXxOnTQf6WuvqpP+1uegnusB5Y7Bf+wDzqVdbN1
EBmkM1fAi9gap3o+1TO1eq+DkhpoBSCNCp4pRscI+wiWvloZeogljZeLPzEpbNdcfriToiTPQ0+p
jiRXYG6iS+JjlF+BFTmoHsh79DogcW8aNrzI7uGhz5ziIadRjp/z0aRgKnEIr31ujGgiSgluznRF
DTwSEidHqfv5Mgj0oaGm6SPVhkYqd0SxuvLF8IMWPPUWo9+qjo+CZ04mkVLcvux/9teGb0NKaa9B
UAtYQsnXk7XmfaWXh+QJ4SNcXHuLVFOht7IB9yEI+Ljuf9iuT3Lqepvs3YPZcuharyZMWzWoTxWV
d8J0swIZ0N+hU6NworPlhzWL3sUszGTE2WPtCGEHl+qjwgOBgDm4OqdC3FiauDSnDgHR7AR/Pt9y
wclhW6G3kqUI64Y8/pgeuuY2fpE3lamsT6tSm0IFKAIPWrtI5WHX1ugTWnSN5Y79+kQX/MmwGOK7
8dm7jr7hM6/xjybvG1WLbzpeSWxtc3qeqvDkNSuQ6oME37ezf3sHQsRgjspDx9FtC8EDLUYRcZ77
o04fUGWDEbNYuZ6Z2FT1PoRWqOI+9OfOPEoco/UUyriGCehvfa5Bj47oeSqgUcMqbK8DnT4qGpxN
H564Taj0vy2X9XNe+IHyyLMeFpiRsZLdZQSE9JnMjXk2DMj4wwYNVC9r4suTZqzdmfGL4XKNeYQj
nrzFXsuk2qCmR5Bp7G0MhDN1AuvgHHYoV7XomKOGMo89hNKJt8jQoDdZ6RVO8+P+nYUE8OGhkb/e
HLxeehasTsS5i8p25mCfPt14EgZRryp1u863ztrlmS/WHuEcU7JWSVSbx/vEjzx3fOJu0DFb6rKi
kL4my5eDZmXDlkOnXeIghJRb7iNN02FmNOsEbSexagBKkMMWRvVeK8QLidjHINe3Xgpx1khIOvBS
XN7eV+GYZT9xbGRLWoz1UardMS0ZWzOD4Qd3yZXoZiBuOVkRkjzc3U4Idj+FfBvrjhoPGR7Ejx6O
jetexxvXY6gbssHkebUDYxbY43emkeg83+dDGtVTN69ffwZ2iaJCGtTUL8MuaPEV7C1DlNRiPa9G
2TYapUkTTY4WgSDb4Xa7QHrgsLv3ZoyUmeLwolGitiagyr3xtbB93RJ+jQbkWYpkOAxNWMZK3+Uo
HKYLIDXWt0jGERkZ8ggliSznFSjzn8GT+7of9/Q6RPJ0fTVXvyh9Ck/e4t0H2NgkCqQ94RpGyrTh
JuSx5Z+jAfec33ekd7i9LeM1iWCk1dSfGkIVyzRnj/Znb2W/5rlLCZQoyRK+EDYLuqNKXnXpTcg0
ig0Om9nVd12t9MaC4IqUm54MklJL1EgggWwm6PbH++oApszuN1fYSiN6BF9vSf6cU88IdKwQIJbZ
bQSZHLcT+hfBtvfAPN+Dg3gxyzD0PWx+iWpf8p7QZ/+hHOh+r/RwOe+wp3+sJ7ECdU034x6sWJjd
g8peflOJeax8o2G6udKwk65AnWh/sazY0J7nyKoxFUmRXp6HF5a2j031cI3XmQv9rH8c9WhhaJ0H
69OV/20Y3CZfkGjsGVDboQIro7dIiLGs7CULZGXh1iVgpMoItF+U+DAz9RuqIDk9S5rQ3YnAUd4m
f3QBvVuYhcd+kOkEtUjSogtvwshyF6VIGGdR8PfA/9yC+MsUxmjsV/iSKlbx8z/zFJmvkFG5Ao3c
CFxs6pOLw9qrV2H0wdzhNRoC3BLy7rEMh09e1YG5IHE7wefh/49pY64ySCJvcRcQpNESNPgkMgH6
rqPevZ7T69sNdQ0I/SZ4ups5klG5GmN/Ex32DCCFsHQ9JvwALjkSN6IKdvCklW4PAF8CV5dCEx/M
3zdlqtTO4ma0w/Ob0/VzvWi5Zh5wwZI62wI/Dos7KKMFv3DESIsUCoQ7ks2vmWCjt4712reJJg7V
G3vdWflxPBqAml/wshwUAoheJ1ZCeLQokol6QYkA7pWXEfRaMgDA/55avRR8RxEW2dgkMU4wHZtv
tvoo6F5QYE97Ng7IJcIxqIsyv5YKg89wHvcHopSCDfDIyQ1JIDoyBv7zVySIf8plaaILO/HI/cFk
W6tDiyT2+m5Mej/GBpu6U9AsH+JMB2w15AUZ6lcES314/EPoUlH1btH8uxxL/NnCusYHzgHi1Tvo
7LSl0wKmRvzXuwyDXpGvTgGaCXjbNScnkqS+gkIPI4JdYNabzURr0LbBEC4Rp2t/ndpofb5C578D
Z5W/Ay6wruTVQElFTwbw3q1Eo50KziogCqIvekpxDltXTwGZDX79V6qiJe13se5cp4aQrimXSN/c
LK2zE+auKOvswF6Kh7ax/rXATTobMeQX49N3kLpElRUPWAP4EmI3Pc/AL0CwtEse5vZproTuPI7g
86K632fjT1fQYzBsuG3SFQ5Lb2vMbevkgGn+5czSm/JAfH7WyN2fh6X+o8sIX227bU9jhzn5b6iZ
xlPK3jsa1O3hmB6PNHkx8SopyLquWjlDt/MtQfjvj6f+BEIf+sBhMl9DA0LY3nXHKPgNVqz7XenR
5PDlL/DAkaR1aV/8055K9uCEnRGrL2YX5v8zVLsloAMq8QYkf/jtya7rkZp0RXbs54ZdTlmNLHr4
joBsB51xC1N97hBd/kf1Nsd++VWqn0qacqsj85S/Sc2byfsd0pV0XBA0jt49fpxcGZv33i6lsp4e
hHbQV0+cTkhjm7y0KWHxDljnmBBqvXJuO/Vo/ZNC/JFVVnelOSR3sHDSJkMVm2JVZRkBNxNSmNGJ
ELJ+MFBZiTinFFLPyIzAjCVwLKnkSnPyOjtw1O9xS7Fm3kRAeFd2+KT36oxMWoytpPH9xdNmkP3q
MHxD6mjnuQ92jQJirlkvDxFt+fP+n/uZOipex7m+gIVMkAh0RKO+kFAmNhIWQ2fjM3LHri4BGVj5
AAaZKm0jL9ga1gfIarylUliv5LFfz+j0BfOzzaEWEnF8lFfeG/Lr3jZkyUmqaaqPDoc2gatJuCbG
sZDpVbM+LBazkrosQ0BimcHpXa2Jvw6vsK0W6hIZCQyimltIP0Nh71x+iccqnsSUggtQUZpvEVbS
u33c81n2hPhA0ii61Qk5BZH0i+NSqYmRbnibFn/boSvxK8FrCQ6pMxu/f440CIYd4zPlq5VEKjue
+0doTX5bFGVsTudSyIbFanV0zi0StfjwvtSDdQP011DcofGR5S2vYs5eeHMSKuqzAgCCmnoj3Y+A
KzGTEuttRYG2F0UspSroQQ3Rz3SjQYyI1QXZGtYbIwmlwVtYv44p75te6Adtb7kH4fqb4UIE6IhJ
vfejSQZWp3Y78xyDAP06vb0qVZL3nyI5QGKQBr1KyOj5fGsMcSL3PMnHd3I/ik/EM1KOSoLNYKOA
JkTbwRXcAiohtQ0KoGeeXAFVUQ0WvfdF2l4XpY+/PcSUQQ0M6sTOBl7ZKHClQG0ez7I2lTjkCJ/M
QB6pyyCP3E+vsM9Gc/nQobxdL7XyCqzKpSU8x/i0XFXpI+eUDYIg49keJ4qRQV30YyqBCAeSoJoL
SB/Tw/pIeJQChAvjP4INL5oTRgzy08POp54i2X2P5B4shEa3i1Ua6Y3REoH3b5Fr6s/o5cGnUCp3
ARzBLfmVbvWvhTB1dLqn6qBN7Uw6UM/vDynbsFz8ATuyQSVW/jsZgloe5nLtVb+0X9KfyOTZwTYD
9kTIgoYZPo98TbzvH/Kp/H3m2oqt2FLoSNlRubnYCUFZWYkyLw+IM7mZhPC+2q3Kq0rjdCBOhpI5
rnNv1XJYSMxnHwpGaD9EZW0kBb8znVYwCMCGWrBrJThoNgo97BCJJ5KmGjHGzfHlUStZsh0vtRfR
bnmS5PVHgxc9LJnzaQVP0PlXEYnCIFIRXn+1fGaK9e5b63HtZe2L1j/AM9BUyBXCHl+iPpm7lEtk
XvRBLrfd6f/Yn/zoG7e+hm7HycxnfrRjGmyaiYa0sqCNCvb/ZRl0SkLikSMC0gcblj1hRR1yplW4
bJTO2uoe8mZropE3ZS1k4C8or8IEdJ4FraIURZdBRqUv7Ct5oxpUpLQ982hIpXlLau0PYNoZ7dFm
Wp7ZKFgkezu/B0de4PdeOf8NmjPt0eseaCdK2UaRUU/Zkly9uxapFrhrl0+nAVfn9fFx5graSjA2
PjJK+9EQUCTC+KUmisC34ucxdJRb1Vt0IRsINFGuxWpVm0xrQn29fvDFr83vRBB/SaROSfUyZC6T
HQiU6E+ffGIBIhkgha+piK8nzX12wHeXOIlReeTd7c4ajml5FdmkwpomVjYAs37eqr5FAQFMJguR
uMqZ83gxGfj9AZ0ukqo/15wkZIxX9jOm3nARg8PcjwrTWhHn9P/rGQc0g4ckYzq5ZXCJVhJYgnSd
rppWeZkZ3BzMSr7CMBLnorUP/dKCn8OSorjotdgqmE888Qz8ld8CWNtJRlPJvY11RJ/lijhoIZdh
jQL8uw7WBWS/QbM7L17p+6rATtJ7ZBDs9ZqD7hf3+SKRHaK6xSo0ymGi3siXi+Epp139i+XsM8uX
oGUFQPSCnLAyi34eoGn7z/UESu2NQPhy8ssYwYpYQVEp6VetNK5amvFf2Xg7TPG6Q3yLy1AN2gyM
RTNsnbIZsZobMowOrUI6eOVo6xw1hWaIuDNyrVprKxTvz3wdmDK2uPKuXt9Nc1NylTEoyb62fOTk
b1BXUm7g44XoCImaUESx+cjEEmcLMKW/xhXQlFAF8YpC4ZvdCljtGeUEV1qJEnBtlPNRGFo7fchg
/JYBa9vebyYb/wrpS/KeElpuAs+e0Sjd1zqAyn5TEBuniqqHVNW4fpUC/HGZDAswyXFFHCaSvKUF
wBb7wo4yPhRMfJVLKAFTdNp74DmFg3a8+FwC+UH3GHJSBo2J/VzmzuOugKlQIK9eXV/uYI2jTw6f
tKn6g+Zk0AE+WV1NqJ7VlsxmpM0CuXTgEiGqOvX56Y7x1NOyPWIJ5C9rRZHoWhaF2NFz4LptE3Dn
iMp/XXJSuYt2PGxh+bb6iTv4oddTANkpJiImXjXpMPznjnLbE8qQp5/W2Irgm9CTD77VLJeKP9Mb
juV9Lt7o5OChoQxfDGlHh8wFDrzhkiuiQlSxGTPnfQ/tpBAU38yZj+emq1XfyY/8pHRWIh9kWw+Y
Tl5FWLW6kRdhQycTa1KHhw/D7pHNJhYOWYfv59VQKfFA9I7E9Vxf3VZgAUGFaX1o0jAq78la3fPN
rtiMdZmuMtWb/mfPcoYUBrly8QeIh98+e4F5Sk1y+FJeXjqTV81j6w1mhx5N5Mru6veVFOq6iDpZ
avBF76cMOCGR2nOwtp/5f5RY03YRNFyhe9sVF+bI+sSTH0JvMWCJO+hHJCLtNE67QDpasO7LH0rn
DS1UXuw6yCOcitBxvqhDrrtqtcaEbMmyEdFofna9uyySar4Mqz0vyCM4xwNX/r/wVGJKhZh3yAzs
9aMq6AQmRWThtlmWTd6ETIZeaeWTqFxjDHrOUGla5pQRrMe6KhOLQ9P47ds2pO4y+u2lWHsoWq67
Ox1EidYtKRUCzyixIaf8Pf09syFbArhB7t35jj7A0zgItWRQvrhw/vwwEXib3vz0p/N2dS1IT2yt
dAoZIXZKWUGsO/T1Ndx24YGMjMYkBZtyYKecOfbTsUmU0Mq7ivwFQ/Uvft45DQG94VO9sUvIBrTv
OJUvDqh/AjiPqR22SArQ2ubKhhVlMVdQNXQh6I3Ckv6DwwlInWPclnUsH9okT6qI0oENbFMWuqrA
9kSOtg6Keh2QqszhLFYwZbQXkzkv79u/RA1ND7FimIvs3aOKi6dgyIJoTtiOB0TIVCtq0BJA9cxr
9hO/OdfnMxLl4lC1N+BOYh74CutSwpEcaxIzLUcSgCTQvTUOH8rqU50PcCtbRF2eWKCPKa7aF2VM
wrhZxwpE6m1Cch3QCsOkR9q0hJdKUQmGFrJkoU6LA3Ga56r9PtsRiMzq4aISbkp6qkdvYJ4+r5Rz
xTKibe9KPOxx77oUtm/mkigZtid79uyUlk2MYpPm0Pap/rPOmYfgrOOIT0MviXXHKrW+zJkEF16J
snGUFIgDuSxqjdYYVRVOmigp+HHC06zVHauvztTCYfB/0Oj02pO8C6/Msqtd3Tf4oHwnBhDtfGro
oioR1nQir0jGrb8UtTizCNjqEKo1uH+ETwpb4wfyIu9BVW3jBS1ufRG03qxpdym1s+AA1zxsk5Ct
5PLATi7vy6gEYbdoieGuwmNjCzoq+PtnTSpp+OxtwTYChKX8NJl2/gUDEPpwv1Zr4zQvOiP8fIHO
DmNo+t0ADxRalKFxmJDfP4zPjtw3B02GcB/AXNGBUD1HxDuyu6hurKAbtW+UFiMIri582oujHPpN
gkTb7h/qz5uwkF5BgtRCyZ4myY7l0wHSBSdcOXFeaS5O50KdDwkcYi2sjZKMBWYKdAz34pOJuiA5
YyDTXD1Y/9WT8Ws22aNB6Djdo7AKygbPBnXPsgTadrBKeFBnCUSaaPIgIswV7aK6oCBgSHiGEBxv
5MdjN6ftdhW96XlZ0UfjvnTr40/p63HJoCZPA4AeL6Gor/lE7f9Sc/dgj+x+PIFqphIHnvEfVUfx
SrXE3Y3WzNgrgI1rnwqK03xVGcglb/ygROqjHrCSLRXk6Mw53mq3eiK9TblUKA75TnDGn7G1niE9
MgAP4/EUNXR559jj9GHhksFr9e6xWkOKXRwg6ttZnqYlbI7WOweAcqQkB1QDTLiwBi6QcLeZ3Iyg
gYpGW2A7zK7mrycJ9czdRO5PvVC15Tf8Ds9aCRJK+M2MbzPM7Q7fdXlRkxKAoVnxohYP/INCpenC
k9sLJMQ2vAyCgj/RYXayhGk7++zcm3oAnnwD9IyGtgSNrsefRjCrMWWzzdONqZ9TATmX/aYeQcxw
NdF4A+jz5tfM82HdYwU16lfU+p1Bk2Oljd3gcgvj/7LCJXve6NsiKGMYHRuo5nVEOUlnjv/eHC5p
BUOmksSoOGWLyNwCUPwM5ndbjvJki9jb4E0VsiYMx8l9ADfBg49EhADEN4Z9zp3B+JWB7kTJEgqU
f4FpzOuIngzTbxyNtMI8nTuZbRgMbRNxCxkn8yCevGiICxUCqW9jmBbTD70wKe2ti7EScHZfgc+Q
WGsrDa3ZX7awo0x56mTYkhG2BlouUeMxowxjo27ompr11Vtwcau0qcJfBFTbq6/cSU7QBcg++Sto
uPcjlW3N7JT0Lkqit3cU0Tl2DFzvNrPAZp+RzbT0JP9mitFAtchXPbEfY+naFXTocSVqfmABD1k0
o2E4f4qpuVU+oQf6BXYrYkCmoU25MR7qZAMG1FI/lRE1wc82zORfKAYJ348F1ZdKKH20H+ey4HCR
fFJW8IH6updTAwB9D/vOYEkNBzSYcOdOWvsHqKhdR2o0BFHwhhY41VchKKNqNFpAl9WK5Nd4R5QH
SGygdmk7r0h8eRLeZM+EXZ66jZJzHaSRFXDSQqMVDja6pYe44u1EQTG1gana1wxl76FEGNSsKbaD
pNug2Gox+oBJt0XS83Xwx1dcmwEBMyZSYNxljYrBAY4WDBNMNHyYInMAAdq2azSxRdj7EKlGz8FA
RqlCNvwXPIM7UcpgKbgwsDfsVKYuLjjZOuxxM1Oa58F26FMx4NXNBMl46uYsbRHnENSxUcNo+hBo
I4VBCDWG7YqhYELyVz7jiGKk1V96vEK3QzpwryrC7L1Gq/PRV6MPOkPGHHWDdKHiee7OJFdPzHb8
1YFzqxQLgYwHGEN3wg3Lxqlex7R8MG+X3DkOaAbzKrYDhhwSYZKmt/UFYHg8DLYP5ETu2ltLj74H
yJiyuUQpFcGZXfsxNOk08ywWgh/ClEdbh1rmmYxjBPbz62PILjn0RDnCwOGMGjr1rZ6ij3uZ87WG
glU+teQGQryV0fGyDTnfC9LyMDdEcbpEiidG9zOx4iEW4eTB1U3oqIsthxJHavvZfy6nw24WnyQM
j/QPyHVxTXFqrd81bqq7F19T86xAIK+Vw5ajbGdUaYZvVuqjE1OVcMcuImqPTM6QkWu3HPZxemPp
Pm2BZftU/FgZeRBhauOVoEmqfDkexqKy/4Q8GKTNT6OH5uYAHw1QgfM/QD2Tw6M4D03kdQY41xFo
2bW20uq62sp1+6T4synywiVSM2MLxNsras8u4whFPML8kvWG1BJ5ldc/ADcDB9Ae6Kl/lWnJbkOA
SxbCnOxrDVfWLYirP7TAlTo6/l849QIgj8P4I8e0Mlo53ajnodc5C+py8nZXQSjL0ChwTPHex8MC
0POIOpKEI+QI95/yCx0SvX0uDupw3x5Lh0g2vCzsvvAyEXhCVL0SjIHym5unDAnRbyGEvXnPP+Oc
JHOP2244AkfEfNK4aVhoDWm6dKcavoM8ENsLstxG1FZaY89lYExoM10JqT/sR5TXm6QDa+uVLwwe
ygMjzBw6uVgKJVqDaCX++A7Zrc5e6+6whxQYL0zJwkxoD176tKDiAwsWWIaTtaSwkE4IA0ub8QTY
1quUp1otNPRRjLgE1/w8ErIk61oVYGB/fgGXmDdj639nhILCkKcCwbiU+zlnJIuryedDSHODhwrr
5+KuZCtClZq3n/8/LLrTfgRh4bJglMaeQJYyLb4S5aXae6T44C9H0fM0+tr/kFeSfTd1cKRIAQLM
2bS5NoehBInfrPkdQF+Y5q3xv6Egm4fdwtR7/MuXDAsvTs9k2Qhe2AWFe+QVWlsXLsRhm14X/QgJ
1OMgOlVqCFXulRzQFyaSP1dDQ2ZQVEB98oiKkOFoZds285fWG9Y3xNQ3OAu57sA6lmUx1CcxpdtI
y4biI64Fplw05PnA40Kg1uHihoj4v8avy7eff9JL/p/TWM5caIbsx1O1j4Zz+TEW361Htkdmn6nt
8cE8EZ6LOuSD1KJgcr9mr73UEea5juU3FyGE6OyG+K63Q61xOZVd1BGz7v1I4JYAnjawLfEQWXLR
P+3Dmw7zWTYsmkjLkuTx9VcvEoeEs54qJvs+pobA01DIHVT8mkOy+MSfR2bxssIv6e47j1VyHL3V
TeiSE1MhjMVrFq3xUOhce9CkV6l4KdSdur9OC/W1kxdO4v67KjNeR39cb3lxbaNMtBggvRiqhXQ4
+Qq8DJDrOTkYs90vf97XeG0lOiTUJX2TE2aF/Hf1JHQ5C7gXZngEthVnncljWsRwP5U9RvQNjCiK
42zLPAbYbR+Mlly7TTiw3/lIViW/FazktmzpuB1BwW9yFHZdy3Hr9Ejogz62wi99/TJ69/c6vvJp
IcOoa9Df1fgXvPY1qjHwffEUwP/HGjswY0qH8ckxyiT7m7yxSqJdf12/OA26FD4VruLq6RU9jY3V
5HHh+T499bfLq03/rzRZ8hm9HaCwJtquyXCFAxlSDoHSby45f1ndNaHZ/I2NbNJjWAh0Hz8cmR/V
mhPHFtpYEKlT38tFlVxWys6ygZ078QOHNr68GsleQ695qHxo0P20N5N1lxjuHltkgP0JAYXzmt+w
dDtNCBFxMurmgw8Y5WgNjUdX1jWuOOdGLevM4AxoPJ6MW+Mf2AKIfkRVC90DTS8q5QF1u2eTu3Jh
DGZI2uHHJ1yLDI1ROVsgyDWX8davoN7O3i5z/piQ4oaV/GG8TFMtWNk2ODM2A+djM/bga3jeVmvN
ZI5Q1RT0MwnVdECWHrsw+owfksMf/x5mtkH68i4eFPbfE36sn/kLz7s6R5SpuYAR09HaZMQi1aZA
qz/+3oJ7Xzn+J9eHampZ+S1hvhECHEDDSJRJ14vKrZXEF5GsO6FYN0bRA4/nxN77vUtCoqIknXX8
sPPsEeBgE3Rw2717GjQZGdKLvGke3rH28RF69DRoBusEkKTuGm+BS3wvgJVzlXUu5cR0FB9v/xey
h3mK7eu9GeX7sxQr5TyrGZRK0qZcSKxWA6cqfgxbb7XoA/jPEv8F5KVXddcoH+OZEwfcsztqd+FV
tTxYgnvKTs3CU+evVKrc1ISrG60ZXtTm1dOU1Jt3W5zAlYoKMIV5Du5IehdS3VLsZFX9g7IGE1g4
zowzRUAFb7hfvJQpVpDnXw2rniQjCYyyH8g07RG7UT3h68gDUwWyi/hioEzdD5nIWwoNzpQaE6CW
3uCYeF6WzpeaRz64eBsaYv2fmdK5qY3hVUCilYjPeCjpuzlVEwPU5s7uNt+Xx5qZl/5dbNB8S/MD
e/RsPWL+z98pUr5c/aBMiJVfDl3D/4EYLVKeX5Fo1pwb0/GbHGXAvbDq6MZGmNmTE1s5AYa0erwF
VgPuQeRqdx1gWDiljvQD4asAkqJf2nlM3wW9Y55dvQMb6lysEAShz2FHotRYqRIMUybqvXbXHb3e
ZIJBSKJ9bL5Ztuk+wjsUJ9aFgzq0rpvKBQYQe6OccXHjI2bL+JXTfNduBCHNvlULC+Pb20YhB0kH
YoWkV2RDuk2TxLtjY5XXSCnyXMk/ETOMuF9lbuGhJ/4z7pg0O8ZiXztrItYagHwAn6COcnIMp4XZ
Kkl2BwlIEgKOrECnjh48vZQraZfj6Gftr78ew7rxS6/0RRT5xH/wVfExaYGn6uynjxG3X41CkGGY
DrT/meoyStTSdU9CgLWIawCqoGgm0KCRN6+moIriwLjhY335n7EckBiqOZbYPLvOdsHv35a7jXpT
wROmY0o8mApXF0RTG57BeK1VSqoKmlw1WuxvtKDPdqS0Pe8UH8RcXkXGmyMooSdIvRTVdBXIzJWL
fzK1kV0YFH8G8ZIWFrTsP8r453UzEUWHiITBv0piY3h4SCJYC+oMIKUaA2ULOd7+roZPYsNCM9X4
5W4u4zRntiAwUhnE9VaxPMhs/eAzrpkqPx3LxKvYtrajN0eeJStJkiWPl/2QjoiqANVuNR8he+vB
iIU798aXGt0QKtETOrAN6EQooWOqWnA9+1J26creShLPdY6hSxeHWLrIAQgPiHP23gAuBvPxRCpt
XTeAwANatI/r881sWBArFxnvWBNj+lAnEbeW8T5CCtn0wSFWjJShb44ipz4lXqRHwhY9ebQ48WrL
DwUowDF9ywvIIzb0TuB9b3uCgLRGsFoICuhhOL1/VgPeIgNN3iDhBm8DA7QnUG8nBgNNvIicC3eC
/HLpSgBQEhoY3hC+ZKRaIz9LwmyeIm2xRdYf7O5+DPxRjBjQG4cPet48DqIHM3u1QWIaP7HQdlRS
bJ+dLNn7UVzixPVhvfjdVV7EBRAdaOR0vRTJzjRjw/fui7MlroQ9FryS3baD5xNn0aQ71J9Mta4t
y0DNB2t0HE+LwdPsPry0/752H6Nmj8d4cYpU3+ZxJRnu+dKGefa6oNtjhtbUj/WqEhYPqdv1Q3fD
hwae+jemN7B9GpEvU9oCklH6NDNBu44FifPkEu9aERkge7imlLwjlo8v880MZpsMgaX/fJzStccE
YQ1s9SJMcJixn1sX10VgOgadtIZAqtgY1lIEG9u6x8CopQqR9NKbAEg16kfERHQCV+PZvf7so79u
R4XmtMXkx6zRj8q43VJeJzL+79PCTK7vkm1Zao7RaU7K4ESkd+OFHuIXRnI+eafaYakxGO2Ol2rc
V79JqlAYyZn9P6dGsdRlDx7YSCY2cZEoJAs73XU9UtNyZldjT8IoW/GBmIY7HIvZ+PsWPhzmZkWh
EclG3/eXNJWDfojQHG9mwpnUAYqfqiVex5J1QL9dWuNpNFLh+sQCDhAjW8hUYUA5D2883kr00LDu
yDWgjy8vkcaPeAnpHAJKz0VyYzqi9Zi7YKGg+B6NADFOgwtpaNv+zuKXBl+eGlBGQvnDt8FyyKWy
g4oz1CBFBSXNh6Jn5+ZZh2jLeuWKp0RCgmmw/HGymtwB3gnhAZQYQ2Dq+YZUFrTjKDWK0q2wbCPN
oBM6xDhvigIFdBEE3p3I+wlj2rqKRztokiLjDbehnu1FUamMddxMQfZPqYp0ztR6rUORsw4mtfnT
9j8slCEag0BsBUg2QlOBuzJNiBO5SlemPcxG5y0K3hj/0e7K01K2aRQQEkXAJzOvIAVvn46OdNSq
pi5hvu2e2AP3uRToBZAgp2eWRYC1EBduIyuo8fWmJPWgqHS2lZ46IwfdSm0dKMHGJqL8wc9LPnIT
RpQ+C1zH1TZTJy722Jd7xnyrPMcyo9I2YGdj7igOx7RlK+ms3RNQCxA/iJ9LrIFyhHAujAnuAUA2
tM1WcRj9Hni9C7CZD9EUlrn9bMUaFnYd6DkWsPVmiS8WYHaBVVLFh/NWWQrNPNXMN9k9Z8g8NWrg
0X105FBTED34YaVBRxN7dFIUyozjncFb8JwfzKYzr70uKjOM8YjSHiJVJs5gmsbZTjhLtSPAcQdq
0yXyA68rzzLoIyKc3fELn7bOXo637S2dO4DbdO5G0MQ9iEVjQlgt0Bp0XYMwN6xsRdCnKejfMg24
oQRye2/RlYEKgxikL3dgHG8zasA263zgePUJp79APup/WdpGFCzSPc4MuGX50u6sWxgzevYAaluN
HQxICTHgPc5++o3/8+xAld/Kr3gcVhDoOZ2I7LAkGImucpean7gc3kMMlj5yxNLWkav8MZPm89Iz
sqZxJawDA4f1JSuB4HoWSq33ludGCnYm8HcpERvG4DTyb8aShw7+wGRvM8Qp8hEbKJ/wBJHYifUQ
+thBA8sBvV0GnnIRJi1eoQPgPzkNCWU4JqW+D3mfvALZ8v7MguAgzHIfGFMniA5xJFK3DltnIQLm
HDGHHgX0tQYf6T9iB+uVdsSCKETgFm8aKiYZbRA3snYNhnpX+SVftfTXidgWj/WpEYF6gcGZMn4N
/yJYnPvb0hmWCovpkf//6DUy/ekSwkEY+FjVZ2aPp0UbmNugODQngtrIZFfD3Np7yYNq97+uswCG
iiDvEfsQolikB23mls187JSRJU3NRN4yLYstFNa/w9D7Iw6pl+Hx4yl/lDYN3X5DuajIJvUQ4BFK
YHB1CEUDetVdJ6BmKtkyD9tr4QOfE+kjk6QVtEtYdw4iUtOmzvKLPF+UeE65Z189pnuAcjrSjbg2
QHVkikrrSYR+pk4MY6P6u+LoBZ6vA0a/9Dp+DH0hIcVDZyqapjhd1pXwEhzBpLweVAkOsz+tuDmR
84HZ5yDiZTGxE+ruXSLwLw7ALNx+GkwaXO1D8DAFq/JUcR107HDmZ5pjdmX2nJ1SBQ1O/GSCHT7L
FNT7CQHAGGeuytL/HljuDKa+ZhmbaFJbmNs8wO7MJiLqk3rjS7tmchf5xHj/fube0dnsq5ZN83/f
Nnqwp1+55dXmjulMWfE67cdsv3khcPEsOb2DvceOmGHMlBzaNM81OM7YoStuGp3EP9wdgteVC/0j
95EnBD1h8yE/poTIMBlvtXXC6EAp0q+s/lIrkSHCfAxx8G3qwz8aEd++YkjVsFp6HZxaNWCl1rgy
pIiV9b0soCmWA0E0zRx/KRhh5EMpQTLtx3jb8pMz/MM9DbNpnYtAzO8/x77MOnfEI7Cot83ynJz2
2fRQLPdSjtk52DjTUFHErSyVRCvoR6qHFNEI7QUqnzYPPMj4VrGzlU/pMT9t51cdg9Ypr1AxQSv6
a5C3JlTXJmkxmpw9SUnHbU5fUfllks3haZ0VUYqvCZvKD7MAvQTdGR25oVJdMw5VswAYQwpIiIwz
EFyOx9dsRLfhGGSCTBoTYPefb31LQ3SrsjM0p8m/yGSnW6Rrby51HgrDLYnVqTFBln2hrQRGxmNg
/K5SIEEWC9vELj8b/KKxMaileHcjHgjCn/0ZGiuPZAWDmIZouipfZD+ou6MZ55CDFn4KRAqpSooc
x5fQyAEN5DbE1MarRum9k2XL6jAVoVE/urK8UsPbtvJSlJ7CIlU7sszRmgWy1JomE9E38lUN4h+p
odfuv5Lxsl0e6zCLA0jrCckJLkcMQF1pUjo43h7B/wucQiszxX0AiFsFh7Cbciyp3GijFlvXdVQv
rHBV/MCY0vUK8DXz6zaw4DI6odWAaXbvsqK0EwH3SWNzi0WLQ+tFyiStu157CyXYYgec2Q4s0pbH
xd2ktCZ+kzHhBPAN8Y9fS/kolUnfBrtZz1k4UIElHq7zjmSvMgUjbvc+FKgI/Kb9tmRR6J7v74il
zFklBGxCAT0iiUgE06FsAipjJPvr2fZj/gHU1QQBVy3g6ziwe1OK69c8IK1snnruiV7H9fhvHX47
SXg/BkY7mp47qyHZL/aUMphZ+ZeNlU4Lpl7Q1e4PpO3hg4gjIVHoqpANBBLvAvCzfX6/0TFgYkSY
kTxz6gZltHzWdS+omxSXVa17cltSkUClX/Ovq6el3/lJ6ZHSfvFX4FnOlkMPTUa6RFV0pbRsMrUP
y/LNGsJ4zNEy5q3PQvMX3wktTlRCrPrLCkZep5LpsuMZVgbKzjIsaANbgVMCVVGQmtjYei2rRMYs
WreSrbAySr6bqQseyQOpBgRkmHmuoaq7HUkZJQyCGTzAXwE/IHfdL++TRscx5DzQ76LqStStI3Mt
9omhwG6O/UDJyCohQ173Fn3c2Sdj0CqCnAsCSETrzkuEYiXMYijpqIpkgl/PlKEisiz4bmtgL/k+
0X/UjbuwXokCUohAc3v0Dt1D65IGUpG0UZL1m7bnmKkmpabYDbzCi7Ttpg1NssisZl+ND4ZJCMRX
uDE1PvLHMzqkoR00O/gu2adYgMHFmTBwBl/p6dLz98KgLImMudh4U4pROEz6f0rcBXWGfvp9S6zJ
hMwk8H3qhFC2WhKAstDsC+k5tSyBKIJfws6Zo5bmkaUkgv4nqBdw7ee+jw501NokBnM+2fkb065n
r0T42txGGpP+ef3Yci+AWdAcHdN1TqLLe8KgLmkFb7fg7Dexr4t7dlO9k2tR3AOaG5Gxclcx6ltV
0GKP+/Ui6em6WO06pMXp86zn00nGXD6YQlgVFroC0Td9xrK25lfN+21Sr+zSBCvxxKQ/I136Ab/7
HNfZnUhZbHBXOc5SeJfNs4DvNeJXMC47pnM/UIL3zYtE5N1oQ0WCSbIasZxezShz0K3iNEqR8FfZ
ZSHvjrTHdJPjXNQ52KzVF8AJLeEUJxa/864Oq5RtfW6WI4hZ4X5wK+MR2OeZxvyNjEoJg0+3Yo1z
1UKTJRM77gGF1+3azOm2vQpEX7uet7c+3Tpob9tWgW0KcmMww3nJa3kxfnbpakJQpq4dV5nGjXcX
a9KpKuAqrgIu2Y6vDttIU7xUZZAkvZxhShlVmj/L6ukxzMk8uqBs1jaibJF0CIO7WPig370FapGN
YcSQKriKdmVRJEISfNca+KslAnej3kW9JV8N1/1mXt/VQeaC68+vRL9ghxwAzj5F4Jx5ja5WXcoi
K7+U4aB2flR+jLZaSs5hquANosNQSH6MhPJFUb8cF6DExKcZny9VMC6dZ1ElwVjppzCYq+VVhCNj
CgXVHPYvGXNNndEBEJtOeAJyR05d+c9nZhWeQt0cO3P8EcCPsC65KjExYk6NfJ7Rfdp+jMpwJ7yJ
CBjuXe+75/6CdSJ3bZh61zKzYj7lvOZsnMW1McBM8PYyIWOA3i6oEDtqh3Ym1RUSYjDmRNdUXrpL
R+/NcEMgprMsUeCfaHu6tbIZCsVvdafGmhlktYVfVQ6ypgsEPbKfW3AXab6CapSo3nuDrrDV47tb
5j6d8UIj3gn7+bMcZpUmoxYc0+IPFS/jzpvJbwd4PNP+QjwEpVwrS2zfqitma62Luag3Fj5mbFnm
SV28S0sjlpEYeHM8bKJAZ7CUQt8ApNntIjtvlLisreKWLFNHjoj6pBT1xqzH6D3ACpA0UYxhtVfo
dItJ9Pk5/+oXkIlqIAQ66867H5sK/hIbj8dED29Y1BEajKRKTo+lnHZXj5ATgvEnQkXM/PYVBhEC
jXJYRHIawme/PD67Zp2305GkkyaBWHbLyOgeANewYTd52XPcNvRpIYCAWcDuQOWPtmX7s/GTBapH
J8lWkJ3ylgGx5/uO8THh4XVaMwey3x6WtxBRZM6dTMAirwaIdh7Ih4HeOTZF2HWZ6tDORj46nsWQ
L9Bgqi/td9u9wnYZUZfnLbEI7hGNqsKuFMwc/GphrmMy304PXSt4N+teJ2ha+DwcKfGsB58VosH3
DK9LXoISqmBJEVn42i/9WF9YQ3MVzxnSmHtyzpfelw/XAXk38p0n5cOQRR0eqWI+YwLzTqgB7Vk1
FBAreH5YZ8zCrJCZv37CxoOPo9vthArY2CpzSBJncnkt76nQc63hs8bWd3hsfwXTpbX/jOXDIpda
Vh00bPk5W7DdASDdYjzVJIYgnoBJIbcJWBBn8kS31gkBKyklkbRZcF7Gq7qgHrTFbZSaFMSEO/Le
DiCeECggj2vMY8xhN9HZhjzMTQ8NitOgd0yqESS1U9xJwhHm+US8PeG87srkwF3jMEevHNWsjotv
0Y3QcaXHxmbfuypqYoZ3xj1iYa8d4wucOi9ujv6xgFsoNPzBVW7UX3RvqH/xqi54JC7DIiKTOC17
B+B1Mf6WQ9nqigK0yRNH/3fgodX+W9fRMhLiBXns1h0MlKB0yscaUggnHc0B7ZKl42U12henr4SL
5jt1pfLxANNvBZ5GTd0maF1fQBzmmIqeHoUzt2p8O98WcFlh2w5Xii1bjg3eHAm7fhNAX44g8L1h
ZTDHwCyjhqTfNWwziLWb5IzvQBc7aB7d4Wfh5LmQoImquvtv5JfM82U3HkehRCXvEN6T2z8h+6Mv
GvffTTT8vVPvSR4suxK9P7zz5jMwU5hg+oLCjJnVKX6xrh3xicfhil5AxGij3A+oytcv0QcbioNz
B1pa+yTPffGdcAILjOg37bfXtEW4km+71tmmUvRLy/wasMVGo++Az+c/87E3Drz5TT9z5/kxUFId
DzRbY+sKrv6wsWRA067vrIi1kIl/y5rkaBal+YuxWfLjFER8pIBbfJGJTTHSIL9DtRGzk7RJJQwY
rdZjf9b4IpPG3uwbX9YXQXeH/5GSLEpq6z2uytn9j9PQXG1/u2anV7XmaDDsADz+kVijyouPI/dY
aogllIaL6Cfzphz18bPZnlS/CxURw1DB7plHc9bqp3kPcOtbiafmGLwgOwWk6FMfLXAmMO4tnAaz
rmUAGNoQGMOW9mDA1eV8eLjW/pRMBupNXSoxLeJnNIVaZHJAxw1WPHzmKh0uE9ehFJ+j/wCnfKlU
1NLBLzHlvDRbksFmFsXhdGjXhmu1ipXw2bgKkvl52b3Yq4XX6dJXziH1lcQuHR6SpMpTLILOySJJ
wqETsSPgqcyKBI5Mi632dOTl8heIjw4vdnFPQf564aQGjgppLxb+e1c6xTqrz9jTjK9kpPbCFT/N
A7Ct0V+SK2ldUlQ40WtGYAnNSx4THcKhGO0KzTYuCm1mqGSDU5ptD2buampxwIdqNOszzwTSqZRp
enGeIMwWZfl0CDQv2G0JGar2mlZA4Ow0s5ELM+0moi2XbCGKNOLzTqXOn9q/V08mlabIcbzKgzhA
QB4iSRPsKyHkG/U+he4N26OUNxSWnj4m3r/TVPbIb7yk7WsOdzcLBDRUmZVh7PPhVmtvOc2dSOBk
9/dDZ9fFBkWbkjaGtdwS2uB0ZP0UiVCIP07xGdVMLOvG2Nrob6YRhBjCvruRzICxVqea72rA+tUU
8VU0ZmxTp4qdYQmw66Cmue8v/le/dPTd6FAJwOaDQYREI+OUy5ecEm8DeZJbyg48F+AO/0BnJcpW
poOmjzWzkyKBNKlWlLUnRPlEF45uAZVBDLJgpSiL6VFIPaJwVJ4YlvZZop8LqFsSuEfaUuhFYI3T
IbV594Qku60b76eBmQqe5YpZhB+ie8SrmBZnWkItVYIu5ttPIuLD/p46TBLlELCrdqwsI5v8SoLY
+EqCiddsQsXFDuq2NtjCinBGFtNjo6RbV+9xnSdPdUgK6cjFnR2uSdAJHgvrKOEb+7GSb3i4L/zn
0VKWIzAeGaZzZqWHIH9jr1n7x99O7gO24qc+XJhlFclB3DNx10TejT9t+6xdGeDNdTXmRZQEGA+t
mIr37eC3l8RjgZSeB5io7hY5q30+T97xS6mgR/Lph+HmHRC2sUOYYDsB8ruHuP03GinAOcYmKUpz
FmklYBIkD4ur9mm/H4hCw2jtO8vHJTWe0t1Vfv35L37WMayBtV8l6rXf1PbwikQQbdUJl+zdT3ry
Ds480YFDdV/Qtz8gjBrNh74wKdxtAgVLa6lXH+Nj97REwV5Gg2ZLcuvKNHj8pn4ssV0wQaNwtgKn
UZyAfuBuZwng411uUJeDLH3ZA0H+Q5s5eXUlXodV9wcRuokGc3F/DVIhy0uG4oQX+paFVSpK6pov
bRkaXIuorHpHxHiNAP++u0LJ/PC00Qaztqg5rVMc1JYIUKuRuaBphhNodzLeE23djhHzn4CHbSmo
4Fy14A+Itx5ja0GHP+UKXRIPzm8oLjJZ9CzyYgiHI1PEyaKSjy+Y3xktJn9RKm7bYWcbtLJH0FmC
ooMUujuVcETsQqjJBRhYPaXIsbMbNvtxEJmaeQpjQaPH/ZHBNHq737TgGiuVpSPGrTQCX+jDAj2D
FUF8GWkMJt+fr8AdvPvmQON3Yvd2RS/vdWd60/OnPO7xEBEJ/Hbi+b6nfuSEn42Bz3aZj8Nmmcct
GF112iPh4aOjTKfabmvd2XzIrmTTLvwV/cJitVQ27uIZkb0Rw34vjPoqRSKj//7J/N14mCSlUc8I
jd8kx/ji3ROCDJi24dpWuzNa6ZceASxIq4vfsLMvfv1CYnIK9a9JLtra4CAxpZo3Xl2Z0efvhBcm
OyYNI0pLq2MwomwQi6qLTz4Z+adpRypQBQ3dVhaWo6H79DdAWsLZfs4itKUqm4pIGP18ttQ0MLeF
WZD2JKyNAwK3tiHRmWU81RNbht/hWTId8HVpM3cFET6jYZ/djm1JD8zRdgXm8ZkYRSdC0D7//4pr
Use8N2OWJfzHvk9iDnb/B0Fq4J4w56IlDnUSN9UzvgB+FPiXZmhpra7apr0K4VhrdqqHSZIEeVsw
/lpC1zCIuHOaZcDKX9B/+7hYWhTUy3CB2gzBGoIWhhwlfppCSgxe0k1yi3ZGjEUQOEo4hwBSFeiA
ACJDThpTfzFz1jmWC0tl+hOPBeIL05k0XZsMaN/zeXHRQqN/TjewAcAAEJR0zYoa1WnzHmwk8Si9
mD7F8UzBSpzaxRueXb3lNqEMfObAy4KSvL23Akulxe4ehgawlASaiEQ0kQwHKEd/K37mHFQepv4F
LZonFe1mxxgrvY6Hw6xcMpr5IldwpkHejzxZ0Jpj0+TGqr7wmrqGUIn4dsvLNdd9vmVa2RIdC9yk
W3SgqSc5Hs7RxOkUFgnk8xq3g6PhvFcuaHKTxIvuSiXS/vuyNYIBSghPecLBING+j6kK66lQ6V+Q
NR/qqC2u/E5N7IN+QSX8c9Qt5gJaI+f+thIVZdylzatR5wCNRN2hHQsTUqEbCHi2Dh69KN+wGXT9
18EWdpFBeHlg/l8GsgkSdt+XRED2HUebo2YZjhV9MNEMhxWN/0MP+vNewhztS3x4JJutlvXC56gX
/CbWS+/S9F8LVyK0EV7fhQJtRgPLyUy9VUOhR+xG7pQ+by1YoO3jGbuhxiNyEmUXxBVDWVcMdADc
Q6Et7tDB8l1n8+2JK6/DzZTZaifLsQZFpJa4MRyYbxIdc4bx8HZPGSifZpG5zAnugYpFKcHFTyXH
Euef9zkNfZl1wQT4wfuBVhIpKwJF6ndjWsviCZ394wPocoAjNjG3pXsCsD2e9VZLWoROl2H8VgR4
C8+akGxYy6ZvSpmv0wgO7dX9+da/dfmoWZ62CCav4ulLSTsnlNGtn/DN5umcNmxYtCSiODdiIk1j
u19M2DPURtowejisBvuIURBbONum/BWiN4gwf+obTiHpYor8jiehIpM1uwhLokur6b0N/UWrmh7x
3c0yScIVca3bUhj5w3FDqrYw5PGoJYrAYUrPPxzx235/1lL5OxztixaR3AjuAQP7Y+XY0BzU6IQW
Vz8VO3NddJZmZvROWdoD7rMUsPxEfuKYjmyYXSccbruHCWykpPDbKUUfVUVR36+TuUGuqiARo16M
QOdkr4DIvBNy2l2vLiHmZhLevG8QMgYSM0UpoyodczzXo2KZZXl3vLkTjNahcsINiuqk8/nFrFB8
tp+k3ZcjMW0lT0BEdsBy8jSWxuUz6fXsRElnLOQPBfyTibYgrpYGxOZLHcCnowLpuBHos5iSu7/X
xip1cr6215NCWfLqwwoNRd02AEpy8jQRu1HGiTzqgD9ikNVV0wMXvllYDPIR/J58a5KtHfvug+uG
Z6rJmqJf3R8cINK6/QpGBBi/yury7pTmcTdpvU4hOMp8GCk6nosCQX/lwTLOx6ph5D/G4WMWArwx
6cl4C6qWZwlutx+bwlMp1C2NBImL0/gICYSu9Z9QviJEvbfiU0llVyh9+7V4Gc8+sgqnTMDOL0fr
qHpPNSDdZUKWQtjpW8NnVhjVqxuuLcPNgk/Qm5xuwPqZH51vfOSImFFHpWO5UhzXUdIEDaYOSjLA
f5bE8AWpe+5Fzc8azteDnfYx1y7+iKxybuhbCtyw+7F2QJKtIjGPVIrdO6Cc38s2LMKfP0uSm8UU
Yy8eedaeEI+3yUP3nxrd+v1rh/VbKGRbuKAT2A0e35EoQm4Carzw+sLy2SV2FZuAvLsJYRrYnCMt
m7xPblBMJqLM4fed+g+YpnI1gcdEZHFbxQ1EmuSpl/KHLF3TB7i1vpIRvl4vGJCX8Nc4BxllC5Fz
99YEsowRH1NTeQb/zRdneBljnYFlkNzgtIurshM4BKCZJ9GlR1LvPHGCiXXqdZp89IceBSKGc6Fn
zGuQP53TxviIJbZF+sJMxOvrbB1kFjqiEZx27LTGfObzIpb3SawyCZewTpuxR91XQaXXqkjvKv7M
t9ttc2n6R92uP39j1J3RY1scG079om4zeboNkOvjGfJvKs9HWnsg1FVHb7Y/BfFy66tJCES6VN3y
OYS5Xkkl6bcTsCjDO0r+wU3BcAG3uy5qr7tjtN2xOwutc41H0bIlZKSrzbte77Yixm+oHB7Mhpv+
2FCBgVYwmtyMVttJCPT07qoEonR5/IC2JoJTbwtla6+0VABPrUNB4pn90eWV/bLzZEm9gF0RX1kn
o5ptopUUPOG8wQRUU6BiB1HO8RoAWJ7A7WMixBx76gX20nkbcZsfTWqI41Cv1WMVVEExF2OfzuKa
rq8VUATpyi7G4PC+KmzRPoFt+E6l4+eemqmLgIfRmAN+K5AcMpjQ10+GJ5lieZAFw1CSOgP6QHE3
zLq4UOheadn6aJqBKrL2klislTgpmCdupoIhIxWQrYJRj4E831bUSxXP1+L5ID1VvzKDykjDUKjs
fiF9nZtYjDW+gvVAICPEub7vFlhdZbR8V2NGad4FHmRMCj9SzdlfYM/6HBeFTOp8cFTES65nN37P
wX2mauy0CULiAKzZV4eMztYNWz33k6tsJ7EW1q3IuZ45dkSQndZ/snPxrnvpjpKc6z/EDwdfcA2W
FDYhbu/C66eXck7lQhjetuSjusUfF4LyuiR4+DgeKeN3XEZBMsP8/Cf5slGPlErD2y7nwyMO8Qsj
vVFtQ2RQy64JwdbK48KYgE+rC9/aYVOdym91AOvjmUKXHD2I/KAIUw19OZrgTZf1UlduCaZmMomk
E2cQQL9+eIEnymtKCnfCPGpbjQEwUHjn2Hz6igJSWunTBE6kIwOgDvlNyYNtBkMPb/joyM2LDpZ1
+lVKHlnyhHUgSj/wFcxggz9U9rerix10Fmf51N6qDmnlLQh6IRriWfnHthPDjnF8ey1vCoWYFjwD
XtRyGb3YSN5WShYjl3RaS8YUIFfZlOpdoDuA81aI2GE778+ITEHS5tinzub309AxJleTvC8UC+v7
ckOvoilBGRokXw8LGJb3ZrT6D5C2+FjO0fXMn3UeJ8phMXA9zk+Z+a5tt8h/sNp4IXIOQISwM005
NFeZ79cqtMJZ+IMGw76+a/bnLtARmxqrS2a22MlDLaGzifdpotrX3EiprScmPre6bk6MUBPYtrgg
CQmk6XnHwB4ocNYHsRGc1z9+qLOlGw6wQsUTXDizXDK65+G0fQbFfp4ecObcZV+qbxhD/aAylObg
fyqheiy7j1vPmX3Zh11paHbtbyljA5xYpvnKbRz5GUQqqWTcBSF1gCahL3ETP/4hrvtWaN7cYxPb
fD1umkE0JFYJZOa+Uw2aTzilZAGpdvC3VgepDvody+ipzTWbY6GH7q03DNE6OxURGpGHv9DGVgNQ
M7pFSbh/iZ/nZP0klpd+miTgN3BYtpCV+ysfTHfrriOTQy1mB/jlfFMJA+WAMqbvOUjm08aB+cF+
NkR7GCCCM69/5EDKJZ851pj80zfebBrsPo0VmgrQdSIuJk38qN0+9h4UHDv3I1f0C8dioYFbw9xY
t6JPJ2cJwHYGtSePjZJ2bFFVt2xMC57oopC+y5Oz5or5U3gbaZ47KmPNCbjkUzx3zrfpbq2jgzqC
JzSunA8ckLP9W0k8Db65xY8Ld7KXyIseFAXFcYFDKB7crxqSAuYWlAksKxaQbtV0wC/33BfTPF+8
cfk7YT2agVzcGo0FR59w08bQ8auVG0kWR8ZnBSgHF5QIZyMPPMHbKEm4ta3Vk63nUk4xhcsbEQwh
3YwzEWe1hkQU56rkzQKAO9+PgML7lcmF70ZBivsSR4b++67TIRfM+DCu6QXoQuK/Cr3roP3VgpSg
m4rm+pUUuSXVT1ErM0vPjnHz1EwmUMsL0Twctz9WYIBsdXs3NmYmPjYcFGuTy3NsUmp/duQyo5N4
PIljMXE34/Rka/fX9Qx+JcvH8puXGgG6Ap8XzojUSwekmUJlf+u7TVfZC2afVEdXni4Dofpjpn5z
nTpvxE/TrmChFkZJpQXi/Xgy4EMyYp3rW3qv7SkUlbTswAcvSaojiwOBU9RUszTnfdzQDnf+Tpwm
6VRFqXaR4KkFPk0pS/AAYlp15ypZNuWGmtXfrlm09Yhl1+Mw/w+ukp4ZeH2ghFhrWoanXXirx5YE
Z71Y+z39Xt3jTOGtl6DBUj5E7qoRi++5jzQ4AG2jkWgYzUzaj0YiBRztv+fNlJzFsiWYTdgV/TsF
ZiVBFaH5mmf0y9573uzNvC2grYj5ZLvTlULyJblsDUnSudok8q/YTBJEKRhmkErRvaX+grizlFdv
A6sYp5iaOVunMbvkRaOFCPaBZ32c174ZjWeJt/2KdAbnctRExpB9Ddd1nEo7ir9FSTsMR3roRzp/
HeE7jtr9xWlaO2TQ9rvPyokvX53ScwJVEMIbSqpfhAFrixJ0PVr5ZhIgsi+T0qFo0PYGmeSH8bHw
uI7TmQYDArIRUFY3GEF3EMWwDJQmTvRnRKWLf1i76ug9WTu88IPi7bRQ2UkprTxbcuSnlQh3tsMD
mcEdFhqOABaS5kKNu7rUTg6/0ZmGjBDYIpWezLu6M8U8zzZmfn/IvM+j2fRf0rTgNOQ2EBN+Ma1p
74EEKWXJoHqb+Op6EXqLX2NLN6MKfcNs4/jWwGLOZTKXUDeWzxsEbyvang+zK3VLs9qqVKxgF51L
Y+BC/1pbg1+D2qKbIUHi2hloYX/GAxiupL8bAYR7xhWcAHGOWZ4u84IvnlcNd2Yx5KfiDF1318EC
DUbz433wg3bV9bwKtqo9A8CpFcTOTV0/+U2ziAKWgmiy93vrB/u80LYT0PbBsqXCXbTAScpFIDNe
Um3t4Aleo6JWoD0z0DyZDEASEu+wqVENvXR37dX0g79b823jJnFIj/LTEkU/sPJ/g7IP7VE22pmj
sFw+BNDGQZVdIBp9J7VOcyRBskFCr51zTU7I17A23pVCKLFT1VycqBs2Oa4KCR0cP/UWXjU3wDyw
Qmzi/BEuO/PPFaWCXHoJqvqVBZrOE0r6/qld/ds4cFUZMTi7/1kGOs68iD+qA79mybNx/neEcard
ANETH4dCs5/mJIM4ewQbZGu39eYU1K0FBJYdzhsme6vK4/3Nf9f0U+U6IoKw3+dNpc4m9NGk6aw0
L0JOGmcjGYqNLSA6o4e+PK+AvWTQh+0Nr+Fpm5HpM/65QVnGDFtSaLHzvd5S2mMnJce5doZqTIwK
nQ/DQq5W2XcHzZOh74zk8yIK3NlQLHvK0hjgvZV002tX0LEDQBhHXLSXQslkS7dA6d2Z4LNxvG8E
MZELa9Ljy4rRqjpFUtJqsnFM4iSy4keROAyjjpyBqpaePagQbWVB01e9k1v5djFXgaANJTyew6i6
Jve6XijLtoUGwLnjkmgWdTzFoPNTPzr/wj1Ir2RKMvyygNkC/nNOXzMsCgZ4AgweCQNDAl6mED2v
dOT/+dRG/IaENytot3AJreiKDIcg85aomuLjgYqb5wnHC6/Td7ttZ3UfYnlBSzc12CfWWKK5/tOS
dJwnbM5ENqI1DplCRZiyO9qrpa5PY5m6sPwtUeJZ1zssutOdXMKOW4bt4wRD21Hys5n3G02/2Wox
qvUgoUm7EaUy35PAMe7I/qB7jsYwinTHZu9ktOdyIvVf4Ncz7puyFXOJaHu0qoxlDo/5brMRDiOP
WZNWcqMZ9hg0SjHR6WhFfACKaUENe1xkxdc1b0ZrZdAJQYDmzeTVz94pTLON5z8LaFMs9Tx9mhmH
KJh1x3nX2puuhrJB2bjvq+R3OC1PSuaim1Y2mC/qm1mZacWHrNdWj2IHq00reDLamrq0wavfbEUf
5QZdk/q4Unet63C+HQO0EKd6T3R4ocWk9BWpYviyPCQGkrZkwBI3PlzoqGfd6XNih0ymTdBgV9B1
QCtg2kOBFR8kn6ipLBBn9xeK8MMcce5Ok3VqZPOs8c/pyd/OLNFd3jzWKCfyIbz6SIZD0Uw41uAh
hdBw/ITNd1zCfDUdeg7bU2XDcU03V3Q/NkWgyD0E0e7W5NN+RN2Vvw/EQxLD2NMsun+6c9+Jz9M/
njGfMhHgYAP2xEDcsF6FwyO+NW7qcbxNj4LIMkwiZTRTf8e2vhKnU6cSPgsd/Spc0uibSMCojDMq
SehXGoimgVsGmrs1G0IdqgGMjvDdE6CiCWzfpbJ+4ftla3W4bTSPf6afEgGE+Pn42Hr01fbt0evP
jfgZXRwIgxI11mLvS7EGHJUf8hvF6SpnvF1jf5NEwe6vW/4GAIenPMaUZiXD5YUh9UlhZjGvfc/s
nY73Mq2ET6CIyCO9wG3GXznJgJR9559cmKsb10sBsPhNwXfngBTeRbWB34XVtBkl6kIU15vxYX7H
TPYH0TFEhFVFZM8h176VPY0hAHbLHAjy7TjkauE+Ud5h/q49EaZZW7vYAH30DcTCTDuEsvrZTVPC
DKXqszCQ9RObWuhGQqJRkjATLpi/qrUlwRQdxob9BtSamO9c+g2W37PoQ5WTok8XuiyajCkGf8Gw
r1CDDVbFM99tkR135jkVZ6aQYCUoj+yA544BgEVdI07bmcjuHhp+EasDTSD/cDu7/yP3B29E2naL
7bUNMelb/CLWcxRGdmNyPxBXNb6tV6yJNVgNxbRanBFgQd3XxGWv1MOiiPf4IVkDbKZ4SKFKcAYq
C7M0fJvxtloLfOET5nghyRTkNnF5+VBTJWArg/8YvufJ7duGuHeDhw0EOl8UKsjUyGkcTv/b2Z8A
eUMxf93biQ6oJCeiCme91lMPxpx18FNYtvSgaBtJjL8lgUAUkOsw/zMlHHqL+1tdQeN3HwSb/8iK
kTSSuz5xvH5nh1BqXWse2TF2L9ifAmPJPmbbVMn4zdWLqfCjy+geVrDTOVZoCVeHLFyWu6gmiN0+
DX9KHJ0/Zz7A/3xmw+3ho3AzAYBckoj9XkKC9wH98fFR4EzfZJzrEnBA3JAhSLhS5l1Xtd11pW2i
W5I9wA2Ub4Ys1WWfJGZ1jggK9FoHJtP22v3Mm4EaHkdDsHsIzw8gvZd8COM+XB5JRyZKHRJolmgu
sWXHttiQxhk+PCjrQa6dAYWy6Wh8CAIwiASbDyAKa/p2BkBgadpeVzgAq3tT6nIm4J7lZRr9fpB0
nE4xojeQDSOM2ucaYV5i7HbrqzqVltXyAgqDuFN2x04jcZMLVp2m9BRKxoFQT/33o8HvtzfBn6FR
Wi7P/g1wisOqX57RcVvmkKxqVAJhYrsZQcdcqQlb6e9j+Bp9by9HOjkUWesU1KmfT84eeBcUHwmf
S/zG4RuQbsNaKkNaT9C2N75xPukVFSD0EXUcN7xHFkMjwPBuSnwvDsrdoM4/H9ubMmgottsw/NgQ
QoBt5OkqgFnbDO0FrijcJ2DbpM2GenwGY7zivtikt+2WoWdNXD+ApE/3hO+EyoZhajrC0BtE5fzG
8AefDOQSC1jY0oD3RsUiYMdwCy0l1sCyNVcstbiorgZO9q52hSNL4v1xQRkq9K5WYyznEGTyqsQB
oz4Jklh3JM/0/3sgXLxULgGp+VdyTRHXZ+6tqg1jsK0Ig382dq0bNlhr400uDoYYqQVJTIVQd9sS
gGhkUktBfcEgr7iWdKJ8aHTXxo+metp4Z4OHijExvTzj8PcoQuZkcu8e8T0VcyjRJY04DjllNOXP
O1A8mxtBdg9tQXTg5X70RtrOlDaJ0q9sWd4Yo/kwjp2bUJ8+pqFw2SNcol0jNHxM3NudrbzlsVSo
XefUbw3ISwNS0Yu0FiPnVXrUCNQ4E5KDxNGpRLM9DaLcv9e3/hHhK3KW+h8h2qA9aECIh3TuEcHx
q4wBns3XtVnuiSN7Fq6G9g+cYkc+lPtTD53P98mooWaS3d0W5hHewj4vMd8YIfp3erEqqSPRXOSE
ouPP6Q9n4q56/H73+Q1tNfNi2y6u9HTRJHSRdjKwTWr3pjFWRu1+SaYJeFi0n+rRD8i5o2tzBhGb
k9kr6pk04UBlJtXyMW8Wc5++W3zyq5XCvL0PYzPY8AOXjUFc/x0+Vump/KmuVJHdHJOucFfugBNh
Dolh0oH7byS9hrgJqg2nwnI6+KvusL1IieDTWva7t2loQEVABYHaiXlpD4hDS3uvFpl2VqSd6ZDa
WCJN9cmBYXVYztRPwtKOEZecDacRoZjgYzmAfWMA0ywx4ke4LhypnKyPPF0Z5yvlrlqz4XKQFTX2
n4LswlN43Qflm38i6gJf0HBC80joi9MdfmtRVNwKQixVlwX9ooR3wnm5CIVhQXutYGBXMBJCGft8
A9f7PBB1tBbxqYfFU0GYBIUv1IP6dnAgz+LujOCDULtWrsXO1p1UsU5i+yC/eG2PQYU29uYLlUu+
juXPExlZw0xWDszmaunrgNm4051ODrC94ziNGjOqQzV99aDwf72rMhxovAxKss3hvq4JLZjGOC4S
Sskv9x0yPhZrtaov3+fynCdVvvFlZNH1laKHLw+aBneKO9JG9YDk3WN0c+zygikRzdox+gzcZxpy
S3zTlZY061us0gMFaOP+ULLXgrziF29jNHDTBWNXeZ+21u3wQuVkm1ENjSwBcutvYLazROMXkv0H
5Bm2PvXu76WlZtTE2c2pdDoLpw+zpakDOp8b1SaGpmeS784w4ug01Y2Z36xbuhhftRtuD3k70yMB
CELuubFMBjkucXLpWtbByMLYizOx+D9Ib4vgnr+NPoN3/Xck0efJOAlJmIQCkGInlg1uu+bzG1YO
htme12fcvG2mX+apThrrHs23dokiyedqFGaFWn4wy8sWjeR0kzU6ShNQrGx8OgyETitdm5G/H9iw
t7CrD1ZXjdqA5I9xPLuhqESEIx5Id6TD3Fk/qv5u+YF7qJOvPEY3mV2QXAatR2e8xu9a6TEIOhlw
bcQ1t3p9IamZa0p7AaCAkRLab4SQlCzYTP7RDdItrYzdRybeITVugm5ls624DwxGPMFNon73Rv8e
emvEmDMvBDYQoyAeV3wCM8cd6yB1H/h0X/oUMh1qEcWKBtiq3akV8wzG39V7xuhG/pNiyUx8XE6c
+uthO+RhEtTBElRO3yVEAK7VUlGEXCuA1qPLlAmZk0XPzE+V6G6eWAx7rqOKo/zFM8sMqKuBBkEj
209BQ8HJS8xQn/aLmSvR+YP+nWMhh1IZvr2mhWBxYHWeDW31zTlPGRGzIfRh/K4TGoOZcxj6ouv4
GHldBEcReJ5A4SM7awG03a+NBqHHJECJDczIgrcWr01G9KtgxymwWfhIENmZdTfnVKmSTSPHYrGi
Ch0YzW7RG5XoBSA1QJ9ofs/g2Nfuut/wKUmqi62UnxhP5NAty0DG3iv7fMJl8xvcxY0IXDG8j17N
FaxvdmPy0D4lMZTvHIvVUiD0Ts6G7id8Z/o8PUFaB897c4iXAkFd2YzFt4JwvzAIei/M2+cuPmw1
PWAn8iAkwMcI9z9eThpj8tPf1MWW4SEWRIfvfkAzLOXSFRnRvilw5DKfZdRX5r5xVdzBeFgujc22
ghJFCqzdq5E77cdht3AqwR/R8X3zK2YVecARr33t85hHn7daSBgxUk/x4PiJDwQofEcgcdHOAcjH
XfIiWgV5i9h7GSWhNtuxa8KiI9kfw3KHZWQh3AIqroanzHkNDVh25VEPNrJ2BPH08R2db4457b4a
1tSH/Y5Yg7jMGSTauGuqkfiynChQxWgeJ520MUggngRWIYDb8/MtYqrGd8HlLe1bf6txlDjEjh+b
wg22dxy12kPEZSLUOetg36ZTbDh8rPYz/8g6cShCtiufRvYMDOJXzEFrTDush8+Uzh64tW40KRWY
XEcpXxw+QBUdLGbNzz5AN8t2nlea0ido3ZgQV4pjZNR9PT9vrAbjhlepFQqEfeikbiR949Pw03PL
P+DcRf7RAzfQ0zPF7dnOjPFIS68jxdPyim87bNeoERCxw7z4q1jLKpGhhukGv+w2RhvzSlNtx4RF
QqreG8ZdPgRfwCJLxdyWQ9fT/PFEwIbGr13eqBQFMaOOMR36cikFE6yI9xW6Q6YthMrnfA+cCCRz
IZ1AHfzjIqn9r9QoPmki5rcK6/uPNSl8bU7U20JolUGjxctmvvMGIuBNkl4iR5QzTxoFDBT4nP6j
Fg81FxyVmjCB5PTTDjfgZyk0OCOReyy8sTeUBw+GKs/OVrjRuM85UfrKJBe54EJSSZDA1UwOJRgU
0dndYazQLwQZOFn049DVboyfS+jM95zT9RWkLfofIhWkBfwaMnAhovrGl21+bVRwe8x7NkpfbyBp
XLDb01DZw+DwCl7sSHxiSuJKNTiufWGYrGP9kgV2xphphA+vkyf07Iii+D8eAlB5CX+iTGzwvisI
ZJdhEx+Nnm2lR+XX1LW/vRw5rPXLzsNOFAFKsT6o5lHQ2v/Z3d/U6fAA9+H6LRE5CMxr62rJYwyE
MO3KUSihuDNR0ew66XC/5EXoXxvdsjG04T69Z0wxX4jM8ZfjsE8XMLDzvIxQVePRz+9B1lJIrfAL
sVlT778yXk1+9hqXDoKPTA2rbkvZmcHi8w2WgVy8nHLmDvJnsTQLSQ5pJajXTsGn5Haq0D6DaFiM
QFvTLgujpiU/uckFdrXwbttS1z687YNGIAHPM2NT6qkkm+XN79NR9fPjhJTfGvniLWw+5t8gGj8I
DPnQeMe4bhIKzv4q4Y6NIBn8m0U1+RQLtjOs2n9BPOdpMG6GRoOciX31FmrbeQVJTy7u3/ceqC4/
0qDu+SlEnZMFObhYFOx/gBQqIyQsF6wbtgs4tVwMs5oxhHs/3qscaIbVpOEJk3VtZKsbn2LsJpUr
440izKf2zFNbYEF6MskMg1Qamy9hnIk2vJiitOUAnG17YWmMTCp/qxYGURfNNFhpil1bgoyLgdJu
j3kVsVPOiCFEdaBh/Q0MLWezHLu3xGaqofRFDEnnjC89GUKU2HctqKLm5ZsggZdS+IQuC6i0AWkf
X0lm4t2RiBoZqAZdVt7D+mXk6ZOUDOlgEXjHPIl4NpPkFqIAn9SfwWA+U5A9KZdndhXaQdqls1dW
ePoXx5RtJkQgnRJCdoblrfVoKHb0Ds2AVRfMicF9fLg73ed8hLgPcb8jsgacBuu4APLuRTG5w1L/
t3Bs2nRDdqrgL7dh7YONhebY2x4Xggvx52TFtubOVE3ToVWCpFiU4In5KkFRZ78LHCmFcHaB7qA4
IsLR5DdCwNIiDcTq2kFlBtHWUhvL7rWZt34HAlTTuw7XU9Pe/D0j3EktHjQ2Gz3O3SRn6WkwHin+
dXiTbL2pAf1oU/Ms+vFm9h1isyDqTut04+WSgQVFdjqlymOLnir1h1NrQ9TNWVnf/OmGCNeYRT2z
SblzhP+8HVp7Fsvx1IE17dNbBUflFbsm6ZgvVNrOpeEbq/aKu3NUcbgNIBpoDRlWxj0p6OTNeM5O
zPWlCwJywsseyXxeVPwfoHV5NKnciHsUulD65KdrMSxSduurm2EZusY2ihU87rh+uE3dOjVKOQsa
TCZNSQyiWPNOttqlJ6lMcAd9wjr3BGW//uGMx+MyvmD35zlKYctxkldjb6EOWaI9e8gDjJMsx9eq
DHW1e45I3ahXAAZnT1CJn7IhAujunxq7zcxlraTLO7qp/y58v6hC70ldziZkDZ/JZquPKeiW40t6
00PaNOXNZ6KotdVHdrv0EI5UyvZbxXIf5oIheaxti5U/C2Rp8Le4y75V8Pf9p7QyjeD8arLvwfu6
72+BEvyp5beuOO38J4XDUfYYPtMGrPjymZacKsaAb11M7l1HZ2MMEuj7XD2Ndvc+Lqih7782WM+6
AXSaW8tKlWhCLHxwrKfJ+1Ep4bcSziEVR9GsBjlC3wH4irbxpgsL2p6RIsu6PvhjAz7AcLj1a1Qh
ZNHmebJSe/9tSESTG62mVmYDP8g3Joqr0Rd98/hk88LsCiaL3Hu7rnFMSNIHNo1OUsuaBXtWZbjH
+RH2B9gPXDgmH6KB/dazgmTcxrTPug0FrIKbkDq7EKNT3H0SSgaaYJQ69f1nDKeXErXO2fK3bsp3
Xzwdheu3+HmoggPed8ZavNSatZtl0GeMjtphgWIycWMIR3u0kwAgmmJniKqTsY/f4SI3JFvCliKB
fZq0ecvWl4SZNNSuFtWdW5nVLr8MndJfF3sfuJmQz2q48a1mjENy4xOtOcBvZlYZ/OMGjlsrDo84
u6K9oCl3nNWzcSHdaTpGMzfhDqi5F8qP03ET1xc3deW79X68EkD1LLq/UnGe5/EKXQp5iNlnqmhy
whYtucBxPAEKBxW1m+YX3cYYwLSMBjJVxc4Hy9OQ3Lgf0b4zCvcxc95e644jRBq4+mAozC6S87Qk
m5KM4hBsPCELSSeuoMEPUwYBMNd07ffzQAmXpjsMH2oCh3FEFbf6Bd9WjjdLyBl8g2rGb0Sfr8cT
se8M9n8SrZ5RkBlgNhHFj5Nj/PtoaONzy25ujb7vuagZy9uW08p2E3TpO/fwjavt021HWiSwzY2x
rXoqpJnp2vToZ02PksTgqh2rrfnNHZVjiBPBQeR4heVwOJetqVpolNYJ47gS3VBVjs6+74BpnZn+
CX64LAlqTlHibuSswo80zjGRNdRnkI9NOUosfMQoMB2uGTn/rK5QFJe9OUE/EJgF+fUlq1XnUlAA
AsabqWlVnHu1ujoxqvABfyWpq8rUG95z8KRR8oTIYXaZ8a2LdijXudAXfS/AobbP/sbLod5zo/34
j8zod+dwvQuvqzkDuc4zs+ypDq9dxi6iQkyDT9l+a0w4zut0E6m3TXhMv2K0A6RASPcKyJ7YDeXy
6YMqmkcc62XVspZUPJZa1PkCH7mse2WZYbsRPJqZCBcr/F+YLtbkiS1TkWOUCpHXsJ6LFlEzlsdg
zWSgsYgtLsoHezwO3Ln9GQPIGKTAIU5lm2oGjevr8JRPDJH2RVEEFRphenu6BOiL2rRhroAmM4gM
hX8+csqZAMkfzFlynhm14EZ/yE83moExcJ+Ba8z9oAXi6jNcOQFryiD8D+9G1hCpYr//yyOcsFJs
O/Fk0qHjO4WS2vqrfiYm4FF6EnuY7Hv8rz+N84ETHEVrOtptL+eN/leYk5r3dpELgs9IZy9JQY8A
W1VQKnp8J3rDV0VvxydXW5lYekCzwjr2y7A3bR+Mc2PDXBkZbQFy4ghZr/wX/oanwz9J7Qj/Fd/U
oYO7/jsFUA+2ZH6R1MP/TxZNS1tul6PQ+OLLoXibHZDmdzWcv85Nn8zImQ2OyQnCVdBp2UfhRNok
3XgFKFizBLuzR8tKPTw+1vHaR4cvd50hbZUpkofIcnUObyoGgQI6QjS3neKmWU4Cv4/kmFGiT6PQ
sNK3J2csnyXhfxO/3m/7ytsnaeNaBdUlD3Au6B8F6muumje6wmIsHrGW5+bULhkjU0/+pJJeoMUG
HMKmxRhi/yAFUuiaMcj4M6DZ4RVdfn8iLhLzvwz2BOz8GzIBmN4+evN6q/1HcN9lhNMn0Hl+MRYR
I/FItMUHJOdS+CBxQcwULl/3mKaL56VCFBDU5Wp1rUPYZxKZDPPhbq2UbRW5I+n4Gbnzt61VYVuy
rW+le9NWs5nh/m6smjXT0iSbqYkWJxJHgpfZnQUcK/Sui428ncaEvPmCE1TyMPggy1nl7Yq/qEsM
rmpUJ0jDxxnxIGoYq+gpKJ2HJhY70GIAH2lWO4+hWRbPFEB1HQJ4cYtS0V+5qPeJn6yYKdl/LMSw
G92r9KTEtgcKfwB07jppeeWw0/ghxljw9kbHPPDZVNqWe0sENxFEEMVlQsOQgNr+Op/Le+XkvYKv
Xsxk79IflVbKcNqJD81kezRqwLkEwSEeYAUITI82+6eZuyQYZcXSXdbmyXMrifXJoZ7twvx7721n
2ZSIVQMffOTzEtqVHkNEphflzS+04AHdic/XgHlShF/OydrBkMzkAKyWMmlMBIG6KVXUBhY+WUOc
WKnpJUEk01qmkXRYnWblDcZf/xh3S7VOE32j9IUMKE0AXgcsbXSzvKylTKv1YkzHwMPi7bZSRALm
nyy3QWLQhuOMZ/MW9ujOB6BWvjzME3J7kg5Xeid7cu97aOpriSD/nTCiFcHlceFE7yTSuxq4HRHM
1vhPMDxTqTRmnYulnGJpFdANYPmGUFUTQYcMKbQdx3a8avNi54D/04VNbjPhlhQO9wqTLGONnvHW
FRudvG1ua8FkR+A3gNNgVLq7ahHoz46sqVN05PvN410yRMcNfr26e+DTNQK1n9npcD44L6J3GMz9
vExAYsB8V0VWu/r3d0XIAhE0Bt+j553GlEFiQAVnN+RNFTu6w5QN14vjaTamKN1v4bOE8WjwBfDg
gUgr7i2Qzp2iTsUIqzYH4U0gS+wvEljDqrgRxbtz0RSdkJDjvEepfGOvB43Oaf0P4siJ0juxoLgr
m7MGrILk2OszGoAWg8e/lWgU35xpVw7RDIK/H6XTItW+WeMaE/2JZk95xAm9/xHaiM8h32cIwPpr
e5QFTvbkcUARDJJIfrXebrHwu8R6EESd+nVbxTDbWWLv8HeCRFdIj7CcvME6aGZgpLJ/UYjKfIyC
CB6qtlOn89IU9Ne9T9YP0bu5BlJiIP+FNPxbkI47lSznQSpn4RGByUyYpRjmPfvUMa1Hw2LdlhCW
tYsAOE6nyi8XLzAp97cVfpV01D4KrtQgOC3bZrGa7yP0R3YILv3apAUxl1wubR0IUEnA51HNeWHh
11nGJkYBjija3PVgkE2rb5dcJMfCU+u0eZgi/r3pfrF/m4C2DZRNPENgpV9PNu20KOzduDE8VzEy
CsmKsCpaGQ8DkV/0QaEsPiiI0T9Ns1wUKyNJCFQJuPgPXfisI2BH+FRLKXkbtfnY6M4IzGqqkmyH
hsbM4srWJkiX46oFIzzVjBMi/dVSxx9Obs/HThYtN0c28Qwz88leK/+RAY6SgxbUHA4OlCGqmqwf
RtEz2bpyB33h2KI7lQu8ZCThIwUtHygKkKeRh71Slhe4R0psRk7o/z6qCtA85v5SzjiMD7QW/bxa
Tv5zXGD6dJ7j9NwZXzmrMm5QI5f7Z6s8cAfKDYRRPaz9GoSqpAKBzh5Zmg0nvnWCDjHE8RTGlbRi
/323I0XQ51OW2e2xE8ML+S/IwM9uih5rTr60JM10UDtZnw18yTBhETnxYuiIqqoiI7Momkz7YXxJ
XCQMGweezjSb2Bjr8URKN0K5Oc82PcQCIt024ZOK6kTx6TAlxxnWyvMnU3ekPHpEPQr+RzzQmE+x
qAlWIhuJtQ9+8+ijmIkyre4OWSAj9uR9PmHivTUG0NAml4npmDUEwKE6WJvENEzYsu5Jiel+Un3s
qsouT0w2s/TnQz69r1+mL0P435EPgnPsiV9DPPSTmmVu6Fdd8BcuECPP+XrgWFnMpIKFaGWb5Y7z
WhfkvOE73o5aDB1RJLSDoCC0LRsroG+WQEzhFcGxGKWrCWWYqYJ4tOnKqBL92EW8tMa+sk/ZxRjP
Su1levHk/unRORJoa0KYsspd295XT6m6DMMW7U1xfukm1CBUWGk7LYAKdbw/0XTxcEcydBn5g7OI
NhFZzM0JLK1nu5ysNPz1tImwmXIZRjq3CRUlgt0cMAv8JZMeQpjXYwBnMkHvMcOhr/XwAa5FmEMY
wdQKEJBRePaK4JEnWkK23IIohV+wFBYw+IxcSbebIrXjFzJG5dChdST4RgkFBWEnU/nA5e7H8QuZ
FxqQY45bUgLgRu8BympyROMN4Wo9c6W/NUJXbYm2ZHiz/zEg8ACpo2v/VQFuXSV+gs+kJXF5O/5M
GIqROooASzN1QGKVbEJs1fn6cRfcdDYftvJvomj2QAMYcam/yyHQ3wpxkuxmEzQ5/DScJsLcgopE
u1ScDuA2ZuLAHDqgoibGfqBv/0M69jvA8f5DUfkiJVx5IKNxiRRXtL6TcfyJpt5hQ3IluyZj43ed
aqUJ6fmlpXbJIALWN4z1kIWAX3cdxrXqvCYUp0qN5kyFzTo1YTrujjCW35NUghZKr4GYnwqYN0TH
DZafGi3il7vOU3o2ODgFsIzBkAqZ44yK0zmJhGpHOPjQUddxvKByMEbI5rXT6qBQhgFXgz0B97fK
43nNU0o32n0uoPIdNiCR504la4o1A3ubSI2MILhskPWYj/A/gDUXFQaAwo9UByOkl/Nay1OqwChd
9p4Ap8fK4iNeCSGa7hfay05Goa900T6ij0YjHlse2XtmeHn6aizyyQFUPxu/aMWBcZe5807LAkZG
9bg1TAnb++Ao0EE4hdEI1qv5m7rM5ICWDItMOZZ2OMoq6+PY2nGnsc/vRUZDKLZlY0LrEaHmLWG0
G0LKHYt5f6WINI3WVuaiLWINfrOJwm0v+5qclaEQUFi0qpyQ1vJ3ClJMwCLQJB9RcnYEQUp19laN
7MoDgmAgnoHhm3X7+YeqRvNVmMsaKEK5ggcu+dvwqSsAyjpeNZPhJ/sTppOSDGjwbEpljX7hfhKG
dIm+xwqT/A6fnTO9P8NV1BzNjPs1KRRKyeXl7xTRvr7CTIJSDGy7ksjd3UHmScKTfOlfN7qNlggT
3FbmbD8vL83QcD8YKH7RR41/sGVj1BT8cRTI5jwpYbdH43Vmwx3HW4Aq7QsVODGZXz79aFN58Vrk
5Tf/k8ct31JfbpNc552PQ5gfQvS/+BfKjelQXYcv6nDqhJrd1McsGnVfv6td9na76v8o1iFzDgVJ
0AYbJSp65y5FgvX3KOccAkn1XeDiy5mHlIYEp8KvaEiNKNG6QDPrWu/JkRhxkyLKQeOav/Ke9idZ
3BQT8fC1A/llZTMtZU+LhCFib5I89zYza0E0WICHqYOOdMBD58Ex40qNL5RUm3phaRDRIEF2/n+p
a7LIeSoN8A9SO7RXBqzRt13YFcTSkq160RG3oQq2fEoelpFdaOWXJNffdR0qScZFjmJIAf4Fn+ey
fTsarseFo9xxnskHMM3Vf+92x1MqE/7z9mPvdJ64K9/0533DYwUXkebGMtJS9HilAvPBEnUTSRwt
haPjbUrkqgeQHemuNIMxVkQcO3r6ubNL6F2D9ZJYHHNTdv9ZsrzctjzUFUMPll8xgUFLl1gM3z/j
+xIG0u6J7hGBgpIluOpq8LyAgHp+JbmbUDiUQDGLa5F132wYhkoiajz5349pLxnrx+MOArgpazp5
UBxjdg5b8qR10HfW/3DhfDKOh7B3Liksh7zRUXFuy4p0ZPG7r6XCk/57gqxeYEPeqBmSI3AXamM5
wotaX9xygpL8jlrZtVG1Wy82nslGYIcq/IVq0+bHU8+/1MUe0JxgUnHxbbLJdIax12jobB+MdtC/
mBIfyH10pU8F4g4/VhzCLK5jtp450e8fRk6SrD5IThDcSb5nX2R8Z0h+H4NDyERlHqbMEK6lNKk1
CBxAs6E+m+zk2iPNJVUZ/0jO3ax85VWcscDYxQv4i847XHxyxuuiJQYqUOEM06nF0QlOtOkVIJBq
ovBhnWPtzVqatXOgRNN5h+xcDuNs+mn5fDLjXYBNGsDobRahRyPffYuVUaH0SlsVfWHz0WUMAHpT
6yCHAg1OA5dQRyNvRPaz9LFV5PBDWwew5mQVK+aqyolpZFrTIHg0JkCgwmdMSGYuxNrPTpsJJAHL
6YNEQkt+8xrkZvQq4ozhRdSdqtzthR/DeKteLzQrBF9Nzn7MK9rpvE1U1ndft9f2FyAXHsZ53nTJ
I+Q2xlsbQPbhmdJyf9tirY8erGuRoNC8eynb55OkFojSoNXjSbiPSQrYOt5x9k4HxgzJQXD40Ozs
p04GKQoC5OmuHzKKc8xrVg4ogXGLYAfYPz1KHP8zAP1I8JF0qpYA2yx1YnHqHLRcGD1/KwtfptkB
gFdFVv3W6A1dsbnH5wawB1UBURlBq1mx2dqRG+mPckAFPQbZGC2X6Z9q6FOpqvujF9TCYoXU76E7
Jjqibo/BMrX7QhL8y4156glE7XuCeXP+L4RwyNs6aPITw6DXfqHf8OHEIgB8iJEP4I9r3UAIo/AW
adsRvkJnK6DQfdE8mZYuiF+MEfNWFfvBf+uzk7pO+1RK+QZz7kUli1yTRaE6Z3HeBaRJ//0LI5+C
7chhp5xGLrcvjzpmCnNjnkSEDcBitkPkDeUhAf6KBODfUxDJhBAvrqIBdwJ+1Zfpb0ZDSBSf2mae
MHFOmwiViyz4ZeguUS8D1PLpkDhGYmAWdVD5rbVbl+D4/NS6T21hXLU1s8pdo3hWuQ5Oy9601f5W
BAqH+9VUPQgKNTYQdW/l0ASDSxVnLhpFP/gmeB+DBqgh/I4IVjoGYRa5eTcNwbl8YnI5he5N5AxE
spB4telq1geVTY6g5fRMykubY5Ac86yVOBD/iaLdhtkioJi7XWj6KbwLzalT9tEfCmVmW8GWrqNe
es4JX4/XsU/0WSTCI6d0sxodJ73Bhk5znDpMNS1GDA4pKRDCqoZHEFRylvl63j+atM7fB7VyVU+3
X2BsWWHpb3IhM4dyTZ6d3k0uf2bnHJxhtA8U8sDsKEwxqag+0qqUmOmBOT+lr56CDk6wc3AJvbJM
VVuoj6/vpZD9KApF+qh5WJAsZL24YtaY+zJ/QRf7J+V7tKD6yRF4BwR3471KsAlWOEjfRKOmIhql
N8MEDWNDRQcMm53dgnlRF2lQl1ZyzW6cwT06/HTs+SZ9YkYSv/nKpVmRE4ZdBSCWM7j3QNSKNE2V
F1+l6avZgXbsZhKf6pdlY5ro7o00jJZmI5Kk9pVZkU/+lUMH/EHh9ZvLPuQFavh1rgqHNkakox8o
L22lxmY40rwsAaBgKYMuLMgfIQ5ZEvOz0E5A7xLaXxqNy1Za6BWYyay1ImC7gfjSaf9I4/I4lUvL
4rgJssbNnQF6CkbjmSQ2y9/KlIVJ4jLw1Gf3RE3eUekJ9svpc0JbTIfUTPp2/nhQSdj6QKACNo0c
UEufa1lKQB+pJqJw3RF+rQ/HTTXYxCllV1aPrMrG3gWrr5V2eVYn8HCY2FqqFKWtU9cHIbNjd5r+
sy2JkX79ogGq+tI6gjWE8sW8xrx8+6ClCVmyrH/5aMIfEmtSTpiSTUeUaRk0D0jseoMXiBnOeebZ
XjuYeYchqA6YpQmu4pfDuPWHtWu8+2nMyjzt8vH8OZnDrf/B5JPkx6PeG9qQcwKZwC01oy1girEr
l9iA5a/5yjkFQ/iSSBVqYw4MibUMPCrbQstEhI0ZVvhOVbkeKkXG3VBe1bY3qnBhfjIGFNOJzwtZ
/jSj97eubLpEIKVwjI//NWVb/3YX81PxLuVfYuzxOIcR4TF/CBpC32RE2oWREb5waeICY/sXMv04
uLXupXBe1Ra3bqFEL8k7PLpuI6ylCCMzmx8yEW0MgY54BA6Mm9ALlsiskeznNhaeF8+vFlgPHlP9
7zwpAfB7xb7jkB/KOYwvPq2rSQyysCijzSyC1bPvo3U1smZfQuOqeMEDrlgfaHhMDQCvvU59Nl/X
qR1FnAUe/nD99/esFxa9GpXlL71OIlabH+JZsVuS6EiTVR83g83dfFizFTOrPvBH29puAj9FYoLk
6OnEMNuAPuZUR5Z6Qn4Ar+eHZGF8iqe9WQIGo1eo6opfCDWB0XR1vgEzqfVndMrpzm2wjf8l3o7H
yLG96WPahnpO38xfJyyCa9Qn/zxLUzIo39IuPu6CTtAKi0AKe8zOvUMpIZa2i/jHS1qGEwEo45cG
rwEKxCAJDl144bXsj/4QZm/1bjNa4A+bNU8PQlMXQd6USomI96CdEBl+WmkSaidJIbCF1TJ+oYjF
NvmH0Dl1Xu0BGbMd3Ta5i6s4Lp8zjNKzoqSEFn2WQiN4DbS3CUCBGGtHtJ+x3EQw5uRKm9Xtwo83
t2w21GFh2Nsv1tbBPoagBB7p2DAtSImU7QHrTgY4UvVzL0iQH+/4h/5K/SaRoSG3JIhahyGK9iFT
DZ2dHTKqRjFg6oCGXNEzEQvBcP4YKtQIl+brAMbZ6c+H+fJUZNwsnMGGuSDyIekS9YrmTaHrVKnC
Cj4GmwaTDR2x/a0QEjO/9xDV6Fd/2Xsb74wW9b11SBUBQPjrA3Uhl937eFW7oV4Fhjd97S5IONYB
IfD+cqr1nhha6ACz60Agpybm+IPe/Ik4cTnz5nhK9IYDzDMa3vW2JeslN4yGETdlFVqPeT8aQLAs
Q7C8Ua3HQIhSaJTQ4jNoPqq8IPpgoZZFWmiCtYOAFm4a13WMf49gyRlfUkb1Ff748vn1lAuKdV3r
+dUdCLfOniA3bqHM1tnLR/KnfeyUKde+rdi41i1qTy1+gI7AbDnHtWqQPrQ9aZ4PQ9u95J8YAV4l
Hz1EU6JVYULnqSzbZd3cnTMbgyglPMpWkRbVFOIaxgbKk5sv/Cs6QqaBTTS6xUZzRx7OUk3A4FcS
X66ycCwd/Mnk+4wZI0Q/Vphs1UNqWD20HNFTA6ZnR+P6upsEmnm26OHSMzUwI3T1Lq5ojyP/O0Fy
3SMLCqDdBS4+Mj6/nvJcjtcsI94m71Zai0bDa1WPgDqIjZN6z/h63dfOd8nZtV2BXb5jaF7m3UJ0
P2/h2gGbEiiQ/23DuW28RPG2C9Z5gsELcWOsTIju4NrfLRqsHvyTlnAXP528YzBv2cCb//wDClhu
Woj0TXliJUnXhL6NeIlJDsjrB6of7waNFqxrLqxOpT5OY1n5gLEKlLV/NEmj/0MGIVVFl1esOlOG
IClBBad/4HwA4n55deR5daiHH/Nd4iCR5/zwbUAU3BvPmPZmE3nyWO7SKU3WRcGUZ4p+3zgKA4gm
1gkGWdpC3mnO08dgOnulfgbj6aluJ2899l7ptUF7T91KGyLLVu37QjHHc0wSbMejG1qv0pZLcxyu
OK2TjIw0xXUrQzHuRI6dO4emTwd0dZnzUj2zZxNpQySskJMviwc8dwhzkVwG6ikkvQrjd13aWgg9
+ZocKMb23KnJQRerMQ4Fq/wVqOkX81VKJGLkhLaBh1JkdI5Yswo8cqQcHCPca6T2emtcKM6QX1Al
pliGg+218uog4uaQu60S+S3MgSfXGMTYA1aDr9m+QEyGjHi8n1zR8OQNM4LCrGqO8gvxVfDaXu5m
COKjaoBC6Fu1AKY4PBV4qkSyjj3eKLpOF49RpmoriNKY4vvJJ5oD7YrXqNQ0wF3obNGMOhDwhiWu
QgZeUCUBgFOnHd1d2RTXpgubWaNmEk/lk96p24UJyCv3/5dM0vIzPS1ViB4jSFzdWqb9h2wy2Srw
krlzMwexFO9B+vo72Omv9cIFR6TlPHBnW9NiuTcYxVn5BUsSZ6QJ80AVn8numxqdNZvTrYLZI+Xf
FH2kz2TQacK8/uMAzkN40P6Yj50JVuyks0FRtfIumAbRpdlyV0vHlWDqSci3wjH3l8Rt6PJ9ZBIS
m7Mj7p8fjH987mExjGd9TgYyA0Hbu+vUFRgO1F4yCWrYmXOXc/ojjf2ihd6kp4Al9O8IRj37H8xH
pWssRBoZVww/yVLRtP/d28/V4J3RB5yI6ZL2ZItZkGOHfnqnSza3C/HWha4Nhiq9lS0KImDmwM9s
z35BUoa3K7tndjpS1L1UJaFsl+pTfvyki22TyS69TaATHc59DLHf8JSXlqs1EoRYBOfgpn61rVmx
XInPRstsBOhlZ4OJ50/jDh5UDV5JSj/IkvKpIkXF3+DzpNiLB97JA0iDz/gXOcuVcwE392IWVAtM
xsb/ILJp9GB2vq2JIOks2RIdhf6CZDTHorueBQu0q3qKTODvcbY9rwHBs2uZg4NycGvcHkDQZt/A
wq8tVZURjWMBFA1w6gDiGQbWqQjAKKJzB3Ok0Iq8WVy118cQBnfM6caQPAzVxj4eHs6fUqkAjr+T
29Bb1+GS6RWOFmoaNb+gKfwBmI0H0K4DWOHgdD/Q7x1uwCatnIxcWxjhnsh5Vkl4AZlR83voPaeR
CVT/0MvZLjQyPS/xx0NLLbThPrVSVE3pclhZqbhoEaPsLrQCW01c5zc14yZZ+Qy1XjXAEXx2Ceq9
IodgfaKA5eeLv3Ptbrv/zgJS1sh070e0TnBb8jz1sOmKxtWNnfFaSZHoN7ww3K8AAuaxumaEWaHl
a1JWDagQoMevihgheQczhuggLc9fDevunx35EN2vgpa1wTiXiq6I56urGvBpwvzNGUlXZLEhablx
+wo+5+MBjNQCw5nA24UTjVafAINe7EDtW8O1yBE0VKtXrBnzpRYejRl/5HloOV5K5wxZZz+091PP
NV1ba30rfgD3sHd0lDnN1czOYxDwaZaw9GwU9pfIuJwFIn2Uesyo1pHO97Z1KC0SwgPUBl684aGY
XTcscb6fCEo4ep9BYrqKRkN5awnmnPHRGUEwU6rn/UPo0IlK+6r2uE1ZLMjd5NhC0H+hiKMERkiL
0f028tc99FNHn52cFqabrbkXs/b0QMzpyVkz9UV8ONy+M5p7ez1QEgx7rJz8sppiqR3v5EJ8swz3
Pm53Xb++0DMLXj4Pl8/uNlQsFLIu96gIgTjKhLQglfXf/2Mpc5HnRTIa/Yh3DVwMLMNJyPCELAmf
scKevEkZdfdCXT43teFe9C0GvyXixOM805BiG0f5cpQvR8lU2FStuBNCc3AOJfeay3EkluouYfy9
XtfvURS3KrZEc4j/hTfzDlsx6I6/V6/CUW7hdGLspBKRhuUfyCkKdByIm3cwFdc/6Ttb8NKBHh7K
SREN0+qcz+pz9XK1JNtMw2gsp6w9fLhAdutheG9JWQj9HWhGubZ+M3qwaOgJ78sdDf4UKczrMX/X
YnJkJlQANgDlQJHy3C50MxUfEOLYR6tCQ/H18L29W25+buZQpTLbifIdMuoymTlqfU0ONxd07zuL
9U438qaMJqDlxxXqzvqJUWtWLvMxAgDCagl3xYy7pQrQrMlLB1l3SmyP/AjLVb7DsQbtAoaBRazI
6GnNlNnqsUXJY/+aOa/Nzah0Dv3XqP5pL2PxI9OlpgEnc+kTXQN5PDMVrD13V87FcKAOjlotObqr
2LcTcz6qxliGFzicDbzsb6CwVBqmuW2B3SNhiyQIPz8IijYrluin0HcOqgs/F+FsHK98Kyaoa1nH
LWlpjkvwAXK1185z/hPJ7F+aoutrNH0g5fUfuOErc1yVIi9lpczaMrWCCFwMlZ+M4Jh7C99aam0K
knjOB9QKHP0nAfUcidwVZHPOJmZMoteJGsVngRz07UGFV1+WnYl8OEqeJ8A5tBi26AHV70iuaUVY
10sax6gm6yr0tG89bJNbot2dJx1sGvcaU0Q6ip5KZoGt7vDYXM5ATVl4QysxlRYLzbekiUZQLP5x
rGypdgyagwGeh8nlTTpYvK99BYwevo0BMZ0B9FkB8mzmp5wGkz7C7ujK7vxYfVfArjIV9Sa7sqP5
kobDiqyx4GQKIXEzQifL+ewiA5nyjKG03e9o09mJ/ANwcIbkCi08oaU1qxY1xlyC0V9GHyrKPqfD
Stt9jh/R5bsLpk504xO5MXyvOKuri7rhchyn/D7tFgmJ1FUys6TFgm+0Ven2drmrT+h0Ymu3A+Cn
p2tkFn2aJIQhB8kyzqvzb9iRp48Rg9yCOzPrjHdhfSATGpyPwCbql37A0JzEWUqJ6IVdHv4VfXvE
a/+85apN+w4vWGBzNOMDHtRqRREoy7vGXvkbhG0aTLAEJ2VhhLRsoWzOrI0OKx2rm91If4BpKD6L
WRMGt3c3Qh8bJN+9jVuITIe8uGw1dhxQHq1pE9uBK2D1Nk3JGgvUE1bQM6eyF0SbMPcRZOool16W
SnisNcw2v6bcTaxgUe6DUVtp97mx3pom0Kw/ffdAMc5IGkH6kBnnkG2Tqv9Zs0U0neYbU0PsgqjF
OqsWLouQKxgDBj38qlp2Zp+u43t3BAxFKKWv278id1Pb/eqhwggkDhFzXAojX1gzCrBwCTtQsBU4
DX8ALmufUsG/maDsoZWOhHWzS5FBBMe39zbuPg7pgSx9UrIsALvPCoE2DyCHukLL7LvWrCfWnKbR
c9N6JB4R0h1rTzBAGNtnB2Xgi1fojNn12rysX8gL+xG4n8jTj+bsLe83lvQ0JQZxGlD/LD4oluTm
dwsopWvW1DPEXAjpAeX48vU6PK9VWwqEk+I0pCXTPw/TxjiDATrZM8bAwlVKnyEts6bd9Y7V0kXV
Y5QCOC1ZnHyKmxwgGb762r0TQZSkOz5Qg/qR1xmzjMbbnPx4ZSHT1V6j2sQn8RUWkdtyMURZ2bHC
GOfeoDykMhDbBom02fNTpRF2x2o1rMx2ncULMG4UaUCxGWRHwXOwE+DBjz26APM0coy/d0TNf7Md
HrDl5bQ7EBB27OcErrLP4kRM0jcI/XTNMDxpFZujrZbIgd8S+8DGC/QEyVtb+pBbw4kY3CZhVTNy
mb9fiMLoygoc/zK8Du2+k49RLwTUBfm57oLcpzZIM0pK97glgaqePrrS3WfwcTCbexjkghLfOTJx
yxW/kOvaD78sOcE47bXasXIre55Il8/ibsc2rXJN4Wxvca8HhHr83AstJYROjD0DMB2M/mdsVXbx
hePNbadLaxPScNOIn4uA0hZkJKN8wIa2pfypEJX3ZfzvH7Gq8J3lFKvLX+YiYbuSyLhcyad9LwM4
DWYUmHYt+KInOwO4rJeThjtrszFzEYB9DOdR6SjGHww784G0dthlwKjHgSHD9or6hzKnvN34k9l7
xIcquJTNYmyS8a89outbIo8hh6Dj8+M3dlTaXMjkeVfCA1RK9WHteKWIHhSSjIEc/LWws+9B8ChL
aqI85HsvFSR2p0Xxx4Qi6BRmaXv9JFSvkYBhGIEBxcvN2YZMnRIM9BZD10E33e26ImpuzH7YaJuT
Go98H1i5OtP9rV8+4J2IjyXPU+jhqLIYk+49tq6uwMI07IxfP2DIqLnjnvL0Jz/R1TWsuXq1kALJ
IhDlqU38Z78ohwPdlQCgUokYJpMIOoPXnEeDWCWyDcCrAvEsg7WwAFH4QHwU/pU9kc4W4rClqKNj
ccL3u8+E051dSf/8kWvlVIUhbKYYJJKOQ8VNoAz1BW16YiQHFMcytsE8+7eRQOvrvlS9qozAViVe
+NfAEBiS/cd7s+Zh/1Obmh1RFiM6WeWMdD6ROEjal6rLL+6HjyU95mu0R7cJh9KsIQ5VDACgL7NA
LmG2Ws77vwfe4JgF+iawsPMOEZRLnuhXG5o1chHZHcJ3fj8jgZXLcPwWsl6t16ka4qyUdFQlwAPJ
8yiGIVMm6cBr7ikG71KT6MhsQHFpNnS/HmH8a1VgFH8YDZ7LRcPqWwfyg+bp8COj/l+5DzAqCs2m
sqMat+LU+Aj7juBKXCLSb1Mnk6DVkJkhh/1QQElM8Dj+9TEOi04dUeRY1x6rUvFXM1GkbqCCGErZ
6KwVFq3bxGkPf8gzOK2Z9gcWjVc1QdNWGuI0j+6VYYpFDBgoEqyktXr1iPUqZ6A85EduQ7XkitjY
uMtT53tTxshcJABC/dpi/j9LAaeXKC5gE74XtaFImV8B9XS5W/anp2G6IcVShHza5+BAmMVfh6lD
hSYlzmVHyjGVlAqidWp9v7ty02ZeC513KAbI0Jw/e8VfBNNnEeCKrzUsxaBRHQ2B/pdq2tQJ9Rpy
So//OPFWhBJJMQjqqC93c6qKF4LXIQ6yaXvYB6dkNEqmivqu+Ogn14RAZdPliTn7Wgk87pcXT93X
hXvZaPOYGi4Fhpzsa7VRivI41KLbkINwxqDGJOfTpk6K7wnwlIs3cy2e9Ll0HxUgneIFxIV1wPB0
Pfl6HJVJ7JxypwXwpIUL+uSxouwKC+wpTOzdA90hCR+chTWXMNfmBkfeY7NXhnTwql/+G4hOKMUl
0cELZSh2BQrP77+GVHgqIeixQlD6LfFQCyEizl3wMhAoxRSRwg+kjp5W7R+AN1Y3uSn5E6bR/Z0h
4AyzB+5ODa1hOhLHUSbAr4PvTcewL7JT3lXedfGvpoaqcHanYFUeXtmrtHsFgTszcR4HSUkQGyV/
9LPD1IlpjwBR/1kxxG1yHGwWKLJSAnrUWqTNATffFeX9+nyemT0CihxGTF+AwKxlHVPZbaBeqM73
sN8tLLj6iGFRFTXM85fWQlO9XhkvZDCN78GHkJBAf3ixAGHkQTG3vPqNDsxPcxj2+70PtWRzlm/m
6rXvOwzCYFb2EK4BPxWV5QTzXHfhGFwdaXxZcA7OKhgko/W81xVEPP7Ks8hzPRKHJ0eK8rMfWvhE
IJrHFd3B0neafkRmgHvTxG/ltb3h/uRSTQ6x8C9iCBpY1/JsU9JGv7/RY7HsgsgScpc/CrCtaQrp
QFzNn7CWoQlI5G8Onusd3jh12vJy03cZSOTvktcscrwYusL6MVLktTri+AnuJPdEX18P7QG9EpOU
YWI95qotE64nbPxD27RzcnsQ1xQgSi8vlk90H8poyGLaygLqt5vJ7xCZ9TMGYxFTv/e0tVzM1BP9
vYSGDhGvZQhAS3k6uEDIyRNhBIrLfFD7+5ssB4VX0RGIXLDoQUEpQSH/UWdoZvsG15Q1Oix0oh+O
APaKTOOvtrxFXRH8BBQRInpiOkqa78Ltc1Ql5D+24TB/m/pwvUjj0o3UiiQ2GUrbAEGgZRWGpRJS
E/+Hfo2abHMrpX3yXCkZG6yF/a5gWW97WJgausfOdrGhcAXqIxpGWxalGxjFFfyfy1yxRTIKdfUR
mj392Hn+Ksvb4IYLR08E8kx5RpQdW8ZpNZTGN+CDBKtBxHq0DghhEU6CSRP+bO6LC22mT97OLtAh
6M1FhCc9+QLk+2y8VXg0WrIE8ENZ1faM4TEPmvwTVyNBrE/LbJvVn/UItKIs6oJJYBoU70hMvsJ8
V0LJqjIcbzHWvaFu22tX7vvCcJRy4NfVV4MiVN21p4cf8FOdCBSkM2S9KVysUO5gAT9XN+M3oBRh
Io9kxnbXQu6K6BVITjW+SyH/9a/GQzZ5LOiUYto5mZKVuSosw8MZvRDo9OMk4jaD7uVRR3XXBswy
aHdQAuDiyvyiKubcxUsrjwhOtnxbQ9Z/64RLR0ohwC1VD+BYLPLHvQ1GabgbikY/d27S9o9IITLl
UMdTwJ7lXqJpATNCBYikHCVz3DJexuUHXRFl5VcTWQHnlsdNwy5MDONzqZ0AZXyP7ggtA5a9mHWM
e17evqe/qt+vKkYh8CAdoT6Lb2sLa79NzU8UanPVMKzX2yeiYdINEHg2XeCVnkdMYX6hXMcyrXMH
+sYPQ31qdqmp1PvkYM39PHFeqSlcGkJ9lDfiGZT91xZqjc4HugSOK8hVDYF26fNSu7GlwX9K8wh3
0jm2k9swLgYarmMR3YwUoDBvtMf0HIOadolZpUtVqbmFaNrkz0yBw+LVkbweCtZXd+qVge3ukH4V
nEyUYgYtC46JUsrvwwXs4bfhZ0KUfX1vHayi8H9XDREvLyFFnGmks2TecKoFqbXzpA9JQoKcT6rS
vU6ZqX90nXF7+PN8CJxsNlDgE5XnNGEjh+d3H1bJfn/G58I5FryPjqiP315Jm5o+N2ldj+L+u33z
BJZa++2YBIPagmqr+/3WpUrapufIsksm3jlRlSQqLf+8ssqKMk5ifwaGDeej6cJdVOHgRK/7KwHd
kbNtaiL3azE7VAXW7XCob0mRIgOL6VywuM3cldgCwe/UNjkmvDzCxDO4fXKBn3OX3dphfFJ3szbs
tUSBfg6gLue/ZynAQGA0z6hPEM1wVLA3f5LGJ9WblwZ3gPiV1iWrCvCigApyq4SJY3zI8TswxhbC
tfqSlALA7lf8bdr+PZtacDuZLiDhs0ObNW1mAOrEepNvuVPcCShxtfEft66eonxJy3JCPf5ZlytS
2xb8ncS9PLrvbWC5Rc4oCaTV6jdx1RwUId+Vm8Ow6gjvDdtPF3ANAp2LDCxiZMUTDlFS81xvsCrg
DXHu1P3RDre9tbTjWsOj4R8FwV4EABk/U1Gh02wQcrfT3FEUMltD4FjcAPMP+urCHp+eWpraQDcH
x6H/1kbClBSjeOHEMMCynEsScF61l2n2M3PGtJDQNcNpriL7xOH27ee7XkdcvBSh1bMKHIj1TjKi
gwWQmdRodrhTWcLNtSlR3Lo8p7eIurLktfIDtu2O4tmThlB7nv9bjpV9BEJRdkPzUDVKn/pcnRG1
6wdGb9vbp7CikWLe8sXhDl96UMDWZeikOtfuqLsUK2SrBe64BNktb7IUp++zEwvH4JaK3vx1dxoD
oiaTCNXe4p0MEWMLRUdFEj34e5cakWdr9Zh3VyGmCezNFHfiKiPuHm/0lE4OSEvd+yGEAu+BrXOf
Nj7J+hsD25RVnxJSQoURm3U/f3Vs0O+VXIikLzCLU/vRbFhpqYT0wL80ijvcjUA2NkK4Ag+7QssW
LG3cO9gK/u03M0jZ1kbBVmom2pqgt//8wQUMOQszD6XLiv27cuTdgpgWgA2iWkJaoP27prF31r/f
1GZehhxAeTitWIn5l/OqYRj+RpTGZ3hwT0NFrE/2ECG1HdXIYvnghF+X1lFRNMzBptErEBm5HU52
ARKPH8Q3DjXaIMpnewQgdyQv3m8Ld3YuLaBk/S7nbd6/daQvxsJWD962j4E8gCPTSNZhVcW7B6ZT
HRx3N3//kjnzSvmos3Ua5xVRuEro3oJ85FQLK35OeuHmtmlnMIUxEq4VK045vAhEvpKk5F3FBaLv
dd/i0oUUxxtzJpPud6M3QPwHToKVcRdTTNn97oYOA+w9RlcF+K5OswbNANEN1v8NY2g5TrJUBByt
uZEcwHFuwFwO7iXwFNU9V+hcpnZmJJT9r/X+cIBksrLaDVdOIWFbNsoRRUhOFO2SG5ST4Cy68iRK
27/eRJW8u5gX9oyuH0qko0nu2n4LPn+WR7M5wdvG3U9JJBm8eQh9PFemeSNYuWMNtL+3sYvhllC0
JMzfdjUWBJ2/JV+NuZC8RJHfNsE2q5xax7mG1sLUAfnIq0Sw8SRJ841l8UDREDD9VLrfOCn4ax+l
cP1xRG0JCoRtsXp119vV5fSorkSyu4sKqG/FHRq7PuCkQxmb2SGzH42Y2rBYaIkSCMEk21lBCCxf
3v7lnY4Gwm40EGpWvmC6AUsAyONuLdqMmfPchlZ3/F20ichXGWmH10/L6+m1MB8RNkGAhwoa9Jxu
W1H3eQUoaQA7dmVGTJMjGoyZwPG9fADH43Nee1L8ddCjyeDiDmy6Nnq9DULnjfDbGw76qOElvpE5
yv7KzhTqKy+6+08S/SpC3t8MieLKbf3CwZIlvaTXfMhXql8R+rHPJg/DbmUKYr6V/fAjjHMznv67
boCEmbLx9Zm+9SrgJxGfqkwJcYvGWKPOd1BybYb6BaxxDJBRqB2LoERLNkc32dzuIx3ax5gzi8N6
teWSt0Xc5d58DTLhupFiRo9xejVYeotQrfJg3JI30ql5ZVGhpCVU2KWf7/gYSdGwjpKze5A4Vxta
P51FA/KPywbk7JqHy54zYNNhUs57l9feEMs21KbUd3zdjWpyuxTjWCxJC/FMDO9hfJpfgwCVptFp
gTchIxQdJ25CO4RvX+ZRkr4UIiNagkb6NJA7InVLpUMfHUd12upnS/mdWHPxw6KjKWHhn/XnGEnl
EXU+Lgjszq8gPzCidpQ+KljxXlnpbLD1LKNl3AezjBCM1I1V6R2kOC+0COna74Ef9FdMwJKVOEYO
3EmopZg7+FdsvXUUsyUEuE+VbtMd2s6bfRQX+yORPujynO4PNetN5q8qpyALopDiGWQI3bRl/Rbg
9uFomg2LhbvIMOYZm4QMOPnrqfzep0ax2GW+x4amjMymZAzijtNDuMqvxKRuN2ujQMqEf+PxxPtb
DVqTq34GtzKy9m0XqIQzxRxLRPP1NB6dlKDX6BOahfjAX6Z4skkT4fxHFGsoXmvWk/rjk8TdVNCi
uX8VqRerpnV7YD/n/F/4hSiKJRpW4xsBK7/mNzEx6pe0YZ56Xgyr0RNa9BDKgvJoN7dLvQlaGFkN
eBEDTTs3lGrQh0A4KzdAjZP12jIgJ9Lnbe9G8T+HO7thQHAXl3e6ewKcDD3VxMzMOLlDMrD21uXb
Kbw0OypcTrwR41+S2++hhW/F1VDqhrT2tZnZyDBgpZfCcJqQvGpTgaxBGKzRyxtMr3x9muAR57X6
1CO1dAFRP59hwqQC4Vu1oYDlwSzT4x6ag1idaIS4Yi1bSHeK4n3ZpKcU8dCAfIoE4zMNY+FHQBRw
MrUqdqxRjxPGN9AIeIcUDKwPq2FjCDuSOD72yW9lNG7jNa4u8Bwi9j17EdOwVtTN5nCcCvJ0avSo
Md2k9AvCT+N/ZxRocUhiscRI1NLxbcSiEgm8lvdfaANnphpm7bBsblc2Ms4KZcNRXZ8N5bYN4scB
/8KEEtcINPPmw14J8F6XkjlEIUBnJB64Lfs8R/K1py0+JBWfyAaJ3t64zK3IxJzhNpXC0OgiodSr
vVjULZj9+kJQdmMI3emp3gzhcE+DFjc0gExdBvMq51ggW3s7cWcSg9PXgOOZM3ZtmLwCDVnc5RaJ
Tdj5DusB4hgdt5TCXGy/f31GomD7gYpoj/PsBBX6MoPElbpKISIVMyt0TM8MME/TgWMaqZpRvYQm
6SgkT/11uwHrZA5VnzN3gKBenwoLsj8SSnllDL7iA1NcwxidQQUlP5RHdWYb1/IvIrrGSEREepSv
z8fUwTAC2g1EU/XEtV7Au7Xs5ehyjBXPdH32j88K4yc+ONCcDeKAlUt8/4U+3pSKU6fN8GP5YML4
Wz1xzM4jtYE/WVcj7GJWlm5ap0eDqJbKLvIkuLSpnfqaAbFbyhqtBeDYiZdneltS4W9GBtNT8bpy
S9RPyM/dwS7+rSkUR5nHYZLMhs2nsqrnDGWWEkU6+kYc+LEN3SDIf8In6aCOU/dy6hLW0Me87zSK
VD43bCkhz05DAACjx7sdo066LDz3Tbn1xDNa6tu+4mNKUp6IYCnedkfiJcJlvopt6f2WVTLVeYsE
fryfh9974yBNQDzWKeLo327PzVvS6J1k15lySskZxTqchULJytCTz3t4afgP+//yIwCWrcbayL67
92kNm61TCjhlJf5ddm+iprAHkpe0k1BmVOGBymHeZ2P6d34tIx/OrUn+2Jz8h2SX1/eW154BXkcA
BcPYRuoukj7AyOdh6ldasgUJexkUG/vI0a+Ye0am43Z3O84YU8/9Ii19mewdek/6tS6oTcWy77tn
Dj0XDv1GsvIVFYUh9ADIysGD0zueNeZyVVIuuAlKFTiHHUTEQEKWp9IcW/gEaF68/Iz2eFUrLcEP
K7PrW7SEl/MtoQ6UxyPSyxm7SE31kw6DEEYcY483Zqhy2h9qu0VDzzG2kE0xhKzsQRjuFQgEUFaQ
9m28KXvHVRuHeG5A2Rxl4Qemt36S2Ucp54Sb5CS5tgEx05ONEJGvxbDuZZQAAwyGp6ME+ljC4glj
hL/a1kMbjLZjeKLEtoB9b56NxkTutg3xMMGb/C3C2xZeoYsQ3Bo++m9KakKXItaVXrxQJbVi7BGw
R/5zF+6rRV7JBC4TbPDibyG8fS0JPkRI1Rod3kh5CKToKHLn65LtjY1UQG2282t/hkX3EnL/TzUB
XigJhsYo6JsmLZhO5VE5OBdxUaKypbpWzY7EBuMWCt0JC9+4TG22Pz+C1lBlCYVzNSJM4GDyvF1F
/qqN1uSZTQdFuvjkR9yn/69tLzqkWySa/WnXgX9ioLDAQ2wJgZ18NobOIjTtn+pYX6NuM9a6QP+j
or8WMmgazmBQk9SRZhXpIWQOiQJY1iisncEAqTY96clh19WWwMvc+tvduh2ghrO2vHMbZdN/eEgl
OB82LHqCFXwdkb9tv8D52bnb5fM/JFyFdR4lunKw7B1QHnjSVbO+0eq9IbClzbG8phTghl7lagbD
Okxho8bF0OexoWG0mxftaZ0DFY3/rw0EUyGxueuPpw/JL1JJJKzD+i5NyyMi6Ebrw1BLGOJ59e7o
jIw/5KVsCPr1F+LT0NoYpZJliLvCFQq88rPMb0fgN9Oe7BOkITIIX/SRchz9ZJqS6RLDFn+l5Vvl
7Gqw+oyOZIGW/5+Rti5Zvad42s351T8KRX1+lFiR7wcHeTg4Cqmaz7Yn4g1rh11JC/Mvl4vaVzhy
GFgc6bGIrjaQFNjqf9+JYCj4TtmvCSybF90qK3IcMSSyMra+UKpj2HCdnsfX/y0FHyZe21g9E5JR
XKA8U35zapo4pK0fzHNPHIvhrb1z8Lcy5w/a7W0la3iLMre3+YHz7o6BgElW+UJBwhYoMAb9pCBH
xbK6C6Yx6aVPSYDUQ+mqowjSjrLzI4sJAM+Ae5knDp/OIZ4jpMaeAXK1fTXBua8rbDilSEFTMO+f
m9NFy/5NaeYg7x9Sfo876qO9fufxThOwBc40pxUoCF6URL1KD9vP2wsTFd9WwlkPPTYe9LHtPbDc
djd7724RoscLW3Ik5WhJuBSnSVAIipLzvwwT60We20sP3at2mF+AL/Fow9Xq/tTL078o1iy13EmY
i7lCaFIyvPDN4GKQ8R+ZI0qjhHx81wDCQU/p/LbKas56yK3ofHiVfq0jBO3QQysnphlivEbf/AtH
ZYX8cz+UfEoWODmLz+8/YO36VgjBOVMOq0MXcJkbwtQOSAy4qDrvdzYY1qfdvTIaY2P8JS8B2RG6
F/zgzGux+pcQ83smS8W/BL+lAn20jny4PYISCrCVPWernf1z5oVebUVBdis9j+JQKM+51vPuzsFz
B4LZ/hZiXs3AUZM9TCAlsMheUvRCYCIeOkltSCJaVntyBQxOgEiO5JJNloXzPIdZ0E5Ws804XmSE
fom0AOv4Xj4arTvDTUopCx2r4f+ZhVsdUo4RMVjpgZ0v3X38/maRYtdD1m80fBBMg4IXf5iWZctQ
1oCF8SCEm64pxggY27VF3aDSpmyJg76wpqffTqpg6v7EBeJQ13bYUkUJK3YYbEdQI3mMyEsXAmNl
q/X4QFbhsFrmF/TscoSVcXOPGURlUqEP+ZIMJbV/aKV5Mi9S7n98APWBPTT9cPizJpEa8ga1b9sz
PhWYWGCJjEVVAa0/i89XqMXrMafLlQ3bE2TPhEy0vcy6F2YPDDksQoQklGc6kn9Rk348sJ7PyGdB
ZHHljY4lo2PX75laJJPUh4og6o2IjmVTURgjCKtuwgprvWsfEFu/rXdWzjuTde2KuBrQyIeV28Iv
oLJEM1FjPZ4MRXrMoCknR5QRmoXi3a8SmCy+v+ZBl042jLSwbWpxrHYNwFp5afVbCbcKbjLvXFYn
Fd8C0noSisMQL7SU9DxbKRZk6pKKzdypNKJTx9to1FbYKupjmniXoO/eIjyIUZ2PK6KSqfujrR5x
3RYqLhWsMcfcZJEVVqwVWbe45z2yT/zNUnTlFI7BY5oLHeUSe8hQq9Qc0vo8WHBxO8ikunzGUidE
sxN7W0w/9CTSx+17WJhIbQ4iK9e/WNbi/NLNE3dRqQW8l6uf3/Jj7fHPwXVbXwt91p8mzagHu2wX
HKjrrPawJHJj4x7wClWWKpyMPA2jHD59Ux31bDdrWoo7ST4MvXvk1DJ4Ipt6G+8mJlbdCeMdNp2a
yHdoFYIx2s+O3PdS9snsaSH0AnjC2APz/asKhyK9Vl34gZpIRNnJz3mtgbcE7+JkF7zITZe+6eSL
1kg8ogGBfjU8XacjYrk6Wgup5Ba7IUcqxoOA3FCO+cyv5K31fZOeW/1JNDPqTzFVWCUjEBnuK2AG
GXd1YaQguwMHfQit+cdK/ixyyLR59+BD9qPDwgnuzuTC4KpJMhCbUl7QS+bh6SqeTkULyVAVLYpg
A2DD932goQcPzeoNy7UVle3aVUkhzaydrXQzujmee7yMH2i5pbXSDbJWi8WJxgQca26RhZVYmfEF
i/dLEhgvjdSzzmHfy8TIyspc0XRMB5uOzXwzTDiswuDNYtJwfbIoCd9VV3JWbLDEcY2aV3C+DYqg
6FTt9BRuy5hk+XIn1tslmzbWZXIc8ithiMa0kTJManA4iGzVD47nk3o4HZaYxMjoF8N5KszLtEie
fsXAtZoeVH8QGdU8P6STe+KGLlVFPJx0+60P5WuZw9E05PMOLilKepjxgPRw1xwyyZE7gQ/WCJUk
lpqZByRLYjd+OBu5RHExGjj2T50oXOhykmY2dXokQEn6cNylv+ILzH9K45i1xr1+raExjBripXpM
YBMJe2/iPBdhCXQ0BnpDkg9oPNWzdK+gFf4XpxGRUWHWKp6HE/ZXa5wjly3vWl4nF9uTiCZUktuw
++JNNHBUDmRbol+xDWl416CMgYFKuoCR9bcVnHbE81DvcEC6VmhggZzFAEu29Ee4BHlA4a5xFSDw
KUXZGYq42sclJqBZDC3wTysFiR5KWVhLC+yS3b4p6wySdu9WxlRCA7iIAafZ9xw2/5wDbFLMKOJW
zuG0XS+CIkp2zNOLp9bNCcVgU2wuJx086y3K4awA+wMyz8zBKXhI37ZyyG53uyUyJi6f53BgiuTK
Q4VSvbn1WtSo9hz1nqqmoydo3lOxSGc2kiygEY6nB9dwi0xyvOpaU+QiAdmpOoh0xqtBThj9yQYN
XAkOq00ynYzqPYQ4+CVnki3xWvQES/w1/bqC3h8/+nKCjQ/HWeNKM89BjHa+j3rTDt1TvW2hST/E
zo+BpOegxSls3M4WlMebL0xFQeRRJLuOXZx4KCe7sHnn+su4njCcb+gIw7LbX1MxyYpiizlciT6E
d4AxTuVoZnjwJAiVkdutSkgnKHXMC1+/pYRsBEM7LxSRIma7zbHKhieFLu2J3ra1wEbqAg5Pi7nq
8YF03nkYJtGkSXzVJwHKxX8f8KtoX8s9dchLS5T2DPNBLYMr9ypbUqlvu91wi/pEJCafOE/mX4bX
LYAY+xN+2Vf7pTu7JPGwssMI3yHZ728H5uLw8gsLm1LbJ2OyJdLM7LPK5ok1ceG9dL+xCjkbc0wz
/ghdMdozYvls5LPyPdNPMqKdj0U70Woyp0Cf3x1d2Kki4Zp4AxKDIXbCC2h/rihMRm7+s/Xotl6h
i7vM2Rvzm1FWGkSwX8p+zMezN4WSi8UgLK2cj79O9pDorJv1dUwATNdyUpCruMWr1c+vE8qFkFGr
2wKMspGxdxwbCEFYa2vbRCePZnt912P6VtowPyHpQkijX9WlWo69/TgMjP20bHKDVvKDESeiBS4k
WJrCn1erWRqlMPlwdn75WrNmFNe2GTyNC/EHnWRPhUFO+0sHExLt+DERRBJoCwnsONDcmV39tb7J
nmLzvYesV01FQJdRJtMin6BBQsYlVyHLg/1YWkjEvssxF9Z708MuQLs3XYl0p/zu4EsQHEylU9Sa
vmtmRZOuQto8PiI7Bd3Y0P5Em201ViPKF7pIBpbmHITGC57IqureX6390d32AMlG1GA/E4SJjiva
desUYgL491DGVEzoMeWN30vJ0rU1ezxX+/QyX/QLquZw3Cp1R++M8bYGdwhTEf9ugwe0P4yjJBmx
UFEiWEE8LvBYLu6Mdsr7S+JzHyFyXxGnBGQReCt75LlwSRm6sUXBuwCBcnkcCxTLpKgTtx7nzJy1
DmEEeMAjk3v7Q1u5eJeOUWNriZjAwTxFdP/1aa5fcMH251m6lBtU/GFumoU6JQ50oXyWpAGNwkEL
Nl4pCNNgqoeZyV/IxG+7EA3G4YmPeovaSKeyXxhRWZE54mO/t6EOgco7qs4Vc1b/W6JPDSFbINoE
L+I1ZCm64O1q+6zVGtb8HD+mQzpWaZGW735gWUC/nqBerYWxNpsxayd78RNLDu3f2U0/t2GVAj9c
Uv+600SGyxlYAbIzAfTIX0/GKthseSUG63/j9Os+6eLSzUqHjqS41eokStaWBrE4D/jkrF8MQ3nG
81njp3u55le2++z4v+jZwB/Wiu57fb+tL6gKZI8E+o/aenjQVlv7JohdwO2izs2Oo8HNWtcCO/vu
heMwgqFU9pHwLfh5NcWFhVf9zkIHLG9xCpaxGJojMFjq4v2XF/sHVIabYz1g4V/sX2V7tLEFateW
iWHUjj1J+XDpkY67aQwO4co401z/3dKE58cyd3N9a5g57S1hQ1ckm65YGIC+J59Iya7pSuA6jZk3
Ko6JyhPDRiTrazNIzhhFu39caKU8RjtZAAT2bdmq6HEryIqZChtfiU/uc+EQVaVAefFWBzd5lL4j
kBMHZWb0C6PK1JvGt05qeTVG55yXtgkvrQDJrEERCiGV7meaBjXjmdOxvPc7sAwEZjURvOnEm145
JTqTtp6BZZB+2OyGCPOSvTV7hqg3yhEC5LFGfj0XB5RVL+9oB8mAhkv4opbSCrC9O3llpDlPKt+p
eeZJ2vAtGhblPsFEf+c2CQ88VXVvGpEAcvOG+tQAcY3vaBlzLywg3F6ryNmKozQ0XydkyqVlQn57
il8rwjBZ9L0rnD17JLpcREPKxcmGgLBd5Hk1Sj//BysgH1r4rHf0JOMx2DpqGe+DJPdtAv14iwoS
i6cKeIBHrZPhILqzoWg8H4phUSJLYupj6fGBPSta+87sUmEs//3FZvooonPz5ZgV5RO2wWnEcImX
euEQ8W/GR9I6Rf/NIPtsH5Xb057dBP5aOTF71jpNZE9uwbfXzTr1kt5WmsYYV6asjSTmF3sL+8Hs
lwwe4NbmuR241fNR4x9VEJjH6gXGf61/gDnihcffl4vP6fahymB1irfxisYq/f0EfcuS7gDdwTKH
lzeWxwh9SS0quUhW/1aYZ556rCRiBvogVbIpi535PKKJs0e8z2x2ZTDhOngMQP3YOCE0xEoUf00i
udt8FoeLvRJ94SjrRMskb0aKnFLVkyYkhlBSfQJQ1N9I3FOgQKHqL2pkYjd4JI1rK+hDdL7Jz1Sc
j32NQQVXhga291Nhqy9K/QQVk54aZC3dJY5MubZgq0QoF6PKAIGMdYlg1yf3+hfyV7WlHo7ZYm3+
39SfC/UVBm8x0OI5u8odAZnA0RWQqRxk/8yZmiAolWvVrJGAgnYvPCaoiVqi5N/V8etm39eSb+Fq
oge4L6vQvE6dKlpKYOlo8PtUMaN7r3G9+9o5WAo1xLBDva8A4kTws1u0nS0pk2kOa9UclrOq8RUn
7IyvWogv73eddZ+yr/pycBAF3Z7ECsyXd4cTSpsSiF/rVTTE8FbXoLf99PjQmQ3ALfS3mXo5o5ld
HEL8SQyfz7YW0fOwHA2qZln2+tVC87GtEFvQfl8qnDJ7oQcOCjoC86e+iEK0+M+o/04irYlJV2no
jZJEjPq7a3m85tHobvicI2ELhPmKdd31jxcXsmCZAbtW30suGLqfgRidWN/b8bcr7wuna1JHwF2c
bkpuFoB78yx5BZhRgY/nEpUnfHPBGpHC44yVx4lHV0PlkRbnt3tepo8Dte2GF52hfvGksmr6y6x9
kAWnJAAjmRn4xCB6bXvwfMhcEErDH9HMZvB/H+R0mbsIpUsRWfuidF3eFEdpmo4FAKI2R0b6V6Xj
NxAfzjiwBnug8z2geHmoc18TwN2g7dDaQo/y4Uc+6+1VeIe02uYKjVRrhCK5fE5R9WXqIZbdPS/+
ae+vJoWK5An6ttq8X/jMXH/cLv8OKCgLQZKr0/9FnjrWaqkSkBCi47efhr4x+zhk93C9PgoOQ6H5
vZ+g5ifHDeI7YFcHKbOMtyIn1mnX6UfpWXj2BKIGOiniVMLfT7Tq9IA82iTa2/ibz1uZm2/qiNuH
B9Jyh7N/eTYQigA4rgYmrQ84fNy9sswJdE65mFWf+Cr+8JeaUxe/dvlzQcc6coaz94FHPJBYB63z
WWtYKHX+yz2gCll+rI2eCguZfKpyMc7HYEmm9tEd/nR+keMWBtdE2fykNXV93/dHasdhwXvwdq2T
8SoFIAXagAdbGdY+4QlBYm4qGvCwnR+N5725+QGCnVJy4WQNOM36SSUoKLh9d0jvAWpZihqp8ZRc
kDjbTR2+pwWD0xiip9iGF7cPk9N1MFbk9guc6/uK9ROc4Gx7MVQt9erm87PEXM3LIpihJMuvJ/GU
zAOmb/VbG62rTM/F7Iyoqa0u0BlbA+4+yhq5jWWTfcm9Ns0BbApWgPvBW//gI5DXbvXWrqKneA1c
l6r6Eutg2/tllRWu9tZGMyY5cWY372USTvvPfm791AkFJPEBpepR28tivoQ+dG3/nkEWDbzPbS9R
/mCDM1aeen8MUg16FbnnVTCtNtgdKLEaGcHxioKHrYlrtoqQm/JoLOhpfipbkPiJp+nSAJCDiCr4
NuSEMQ5njX6lzHNOHu2bnZPzshWvRcv4SCgyTFF1V8t210tuAHo2bjw+LEKKWrwCU2u/TMq/0ff1
6q1oHKd+Br5gKKifiToUYWqaw5iSBxk0QOef3Tg6D7hTYw68A69yrGyV6moAMKVwW1YAddPfCw8b
RCWO5wcAX+Oo/Z1m/jsWPmaSnkx3kse/EfmbPz5kciwcBwcQxvGOPJkr/T3zRSU+CS4JAqF+CVOg
54Jp7yXOHKIRAZMNGPlTKbYAYhEyhUT9eLKqk86RZSix1Rru7qrOG7b09vKE49VRLxBc7EuPWHxQ
MNOlXC5xNLdFdF+NZ4SvSMQGz9xzy8GLWoU19qpIXv+9UNccBWXCuRXEILrdnxII4PEMyofI/3RT
lvvxy2T7VaexcT3lQ52Y7/vJ8EGHXX8JskbN0A+FsOsFWrmxKF4dWOy8Sx85R+4F7kT3T3pRy5e/
6qYmnDJ4KHzNy/qixuCU2tBIurszW16GTSuDGq2+c77O6KXejy6ipRBjdBHhHtR74tJn6h7hnyYF
nEFX5AvCPTLlaLSmP75lm3vREWIA84foHX248DMQfeNLJvfHINDC/KF/FPfhH/vd8RtYlEPPi+OQ
/+ktBqy06MXQcZ5Sf/j5CgdtdiqQjreMOAphKhXESC2iT3dLFMmLM8gCz2urTCZW9lHYBt8mBKVl
RoqIfPxT/gJFWnB07wgg/SoC8iMxdgxl5GQS9bKeFmk0gGcb5dlvTWRdXwXgmg0VKrY7XpuHoUBG
J9VEC6WsHWOKD0uG4HIO4qtevXzRRefhlc9m0PDC/k/hgMikZNwsUyNmAJaxvYae2GuD+qtdbpJh
YVIMdifGnTsO4eI+nyfQKitoWW9IzQx+Lh0HZiUrygc9CdYCTyXjo5rZ2UDsYquYWMzdyOs+7nN7
LQzZUD+e3DRr3495jJ2aD8r0OGEqkFLBTTFU51e826JHbNdTNAlpnX0vNjOSNuKBKfIqZRzQfyyw
T0NbANWLocfSwJnug5CrLokdoKQqnuILQdNg/k8Er33a9LhYygvdxyVsnMOQetFM5V7WqEI2NfQz
eoOPJOSmo1q9pfbiUnR99JrCwFwn8LH2y+MkQvOMtdXH6n5yoaoDejbzWPLfmgoTviLn5jjsbWqV
WKXThQM3gJuKO5K3SQVg9pImgnYRtZuB5LSrysryheGbAXcgqex2PrOM417e+ua1tubIrrn2sKA9
f9ONqOk2qakSolShJh+nTDl1uk+wJE8zyilZew3F3p8iXBART26pYD8PgV9dNGzjP7wp6TCU4LKp
J10gQpldIwphEOt9Y3B4JT3aU/dDnX3HX9A+uP3PZx/ZHj1y5f84wKVHFBCzFrWk/amb19btVN4F
MFyaeeXwxCkfKEXEUAjuoZwUhEQe9knj3oaI/429E76/g2NAuu6nC2Q9N5fg2k8BmpyJJXaEuJvW
dTxgM5e2d0AalbuAhEZYQv8BC/4cuEQiEKmBYr378fNCjKnmNHMVcAtVOOnlWkV8cph4if1HFOJx
7GCztwaStuFewP83KLm+Ka79eqCmLMcnfgfyR28aOfJ/kFAI7ulYv+FzB4Nthmla8KomMGD6ryW8
674+VBnxydrhDeJ/liljryY3EShraugVdWSBOEf3Kk8LjbS0H28sGDTQ/C0yBn+g+13dcR0Efdxf
QnMboZWxS9EZ3rM5y9PiAI9NB+9rfzOPwgcDr/vhuw2o3ooQ6Cr5YYIHFzlqusoq1CIk6dxD7lJG
wnZ6J5S8und567Lgo15pacygR2u91kxtcDCRI196dCpmi4BXSXDVEtz2xSvR/P+ka9PPlE1MYqgw
/bUS1mYQnEqRE4/t+PtESH8g1SIxGLcj73HX7dBqnG+wFAH4peApRI00N7d26dUwTqd7vTI3uULT
DKYQptGruN7y4nYdhG3GNywBkKYbL1zsnIl72sKXxXJ1KZr5KyL2M6242yi2Osgqoq4aaF1xPrTd
5Lvn7RN6XbbLo95TRy2JxxYvQ4LEce7DwpJ3nK9CrpdtW2MeF17JYvq08DjGgjKIWl0bfcnToZdP
dDIk1ehZUsIKxiYo0VFcHCHapCH6dOYUIzfby0TDAsXjpqzCdq+B2wegXh2103bh8i/4fGNscrqL
OU1amJFaSTTY40QeEqRv7HHC/qbFFDpVtdIGra/ID5i6ou1n2TgMQIdDlx89M3zctpMURpG6GnMg
q5vq7QZRAiz78jzflMLcp2m7q3/X2i9ieC1PecK31psspzG4ghOz/sGpSyfpnOfr7KNg4b+Mfy2R
Q0jQJBJTN3wH8UHw5Hcd46LaUcRZcF/8rs+HtXgDd4bEz1002EnbWWPalQUyPf74/tebDHwy0BCq
1M+2VAqkDtElRnEjmDD4uVkwPiefDCmoELY6SGwKtzvWRYwunuObblNQWgbkEGy3pC/4IRaoNl6F
dv7AYcutlOz1IR2ZjNUR81UL6+2+Dmibs+phSH8Y4roDM3Xz3ZJh9Bv4Ea7+YHdNaFIsIO7T2VN6
FnmomHwoxlnIUdBHgRDiqhcRsoSjJjn8+JhuUoBzYv57yqzpyMy8WJfcBO7uOeAeOPVSXfGQEoS0
s4g+7vPPM4hPUwangdbFfwFEWAMGrn79yM0opZOh7EMNUAUjnmqCIvhxNYUQ5L0865nx9LDj8frt
sCUDyCmM0Mj8d3Za8mT7tu3gGFe9iQOukqx1NY3j1vEvh/0Xn4VHFRlQ1hXtNHpii8X7iGThfX4Y
XqvfgSmWdqkC+kMo9O0Wslo7u0alpOJDDc2F1FJyH2O3HUPQYzdhth+ckIDkwbYKhjmWHIEVr3t4
F1x4VoNlROafc0OCLqYAlNwMcF+OFXl+IawS810KqJm/gufxJLfD2bvNoJNt9ZnkY4JljZ18c53r
jbrnjFnEDp8B+wXHq/u1aRUWKX/93cMDlxVVvu98B+sdbAsdh2Z6LdLFNtFYpSMjzsKmS47MOqs5
pPVXqwv0GqdnP1q/uxg/Ke1lR0kpntGVx09appc8GN0/czY37Y4SWOhmcSB9J7pah81IIrEJgtyt
0iLQ3pCunF5ks/FhP6LkZEyaAji471FtG/ZK4AWAyU2nBwk9Tw/BhcrOkL8/n+P6kpAJipdQBgtX
eLv6Cw+XQyBBjKRKN0jXwTcF4wyE7v8stwb9ta4l5IUTKCX+OqjzGzA5rdS8vc/RwglGhKoYMPz2
YsDvgnIFKMMrNouXFoZF6KG5mT/lCD7DXCKxzl0UkzVTn1eCjUTVZ2Sr7pBPkAx2E680Kiz7tCUX
YKeXyGSDuG4MH4BLhkeNuMWgOavZwe6GqAgLJBH+m/brxKoesL0Re73qB40Ra9dW2D9AheIIdV9z
QAJVYAXEiNIeT3U6MJeoDaxWr6q98bNgNN/nEfpoXAS+lS4R7mX1hxxWiQnRF1RWDrankL2ANxLr
8pMoaYy30Hc1sfrVMBQpLBrlcmnnoBPR6iBjxjuZeRO8/il/lSKQjCJAMxJPkxBUHaPORfM4oDVE
SVyI2V87qNxv2JfgF/p/IFSoW6gpVUeB8bZMxPu1VHLZJ7Ms3H5eZzfd80EnZfQarvv3KeTMMpbT
1mwix2KHAepQd7LAYfbmcgSnK0/6TDw1VAxPGU2jTII2/0HwUCxKH4xq2WR5NAhc6HTyOpU4BCNO
VfuDURt8WMlrnpmxsQhZt6OYmcDqeKSt5/UJLv7wJOQjob5j+U0b6ADqrWXsZD7hs4LKmotrwW6k
RVdni4IOa7zAGeIdVxiSfoJU89CISqVvgJugtbFrEvJ9NVXPl5vqWDtKuz2c4vRIhIhmD+Oan3lC
T2/vrXTSWe6X3fepFCr4TiMsscACUU9Myq08mfi4bZMtP0lq+CXIdtNqlMnXp1y887gOd1MFiEwz
LIf3eEYgIFyj6GbLLGqkSRIzHiL08FbFjoXlLHD7eT0UeZ37CSDLyWo9WiZW5LhlXvZQqRtF4Mrv
UX/O8CCwYouMImiNP8yj71qUJKpL4f7zA/P9xdVZRoqgOeezly2LP2RWB8+LmUUvYB22yGBQJjI/
mdxWlXRA/k8lPi3w7iwd2GPaAM1nYVn0AvK5FFLdHFU8xpE1YUUU+7uOv0bpcZDWQv4eBVtumkNQ
kRyfIHdzXGLfskbMKwRyGHgx6vmH4vwAC9r8L3WuR+lATPyoCSkXBtmd7sAMCWuhuKiS9llW1QiR
6TGdPUnKdqe397vQE5Ky9WC3muClGBjC0D8pa5P6ik1DILTQvfhkj+6f6cI7AVYDnwt/RWLIo5il
dbEhFbuExcwOi6x9kAc2Gjo7j3CwqiVtfF6oVwEcWdkgKY+HJQy7Yjan98GWafFtVublvhluDUt+
zAirvAGr8U9jiY5aM8/M7vQJUcfDxsiONj8A0p0UnxBNDsV88iEur0AEhAUFdBmyNtZIuelYAWCx
NTI2F6KNhsQ8kPfb1Rk2caob1BY+T8FlCn5Gaj18+aUXYAMwLDDkCaguYi/cVtisyRoD8+292PF4
pzEHjOGKBBFbb3Q/7pzUSMQ03o1FSJAuL/0O3k3pwD1VzcclgAGdJ390vyjOMgvV2VrCwSBOUGcG
CQIr0JLIAC/IvrGD3sCLhi6uBEJKMHE+4DruxHeKzsFWMifEjbJYaV/qk6iIcRhqso5KXhYeEF3s
5BTNYqpnkEdxLdwdGxV+B2nxgbpHQlDS/Rt1QtZs0gRx4yFUJG2TtZ+F6aiKchhwTeuJzrulLCWk
GdaKAAKbK3g13gX24wJe6Sx0uKgInzOF5uc6irkUrpoB+E40H6KHRkxM1DJwOPcsJZGSSR7tUQGv
w9AnEIqPwG7J6ZvrbnNYgxwnggYp9kanzFydqHRyXTmT5tgmv8ppAyoHmivWkWVudxGBwgxQR9Pp
m5ORyObI88vq6Mc2MVmvr2hXFmMoJIuTmrfezzBZbl644XOh/ZrR7IDfUfgGbrfOib299ZPIDIay
Ebbmxm8l8ExFXoaoH5xaNSMhL9cc08KNe0CnOGm47UwYHTVNg0REdw5kmwfJYSuzhQ7+UiTY6pgd
ZjEL378cVHOgooqhZ/L+OxIi1gD9HEGUOOXwtsoSV1diEiD8sLNyuIHfduBue/39d/sFo1ts3Jek
1gcf4Dw62NACZoiD5B2574kS0iYkOVXMjvsSFPW67Qc0Jt19V9bdIvmUBAN7sqNBRyEIw+fOLWN0
SP5xXkT8MoaUD04J3m6efXhqmm6WSG2WZtEZg/KMdIH5TF5FzzZSDlC2fpKZSsR97FolrBQ0FtCX
D1xrXTrW/Zrg+LKDA977rgPSBj0HojjoOQB1LIhlgt87vJt6Wqd78d4/jKU4/klqENjIqQcqsojw
PVirfHciIqDUCGbqXamjObUTRAjln6SfZrbv74KvjTMNsJHu/4G9o/nH5f518gGP+sC+h+3/xrkc
jXAQSdNNYZoRvDwpDB7IDQ65ISX8UKq8308RPCVzmocxFSn7z1quEyOd9kGfMwPMJprYdk/PVbqq
C/lCgbip+CqIkrBIwnSsxZB7xyrJgvVUEHoToHEuQ78LDnjOJss5xnwE2GLu8LR3lcusvmUstXMs
NmtDi0CODEJRchY/G2E1iwGmHT8834E+s63H8YKTM/918CHgQ0bkVWI5pAw59F+m0DdmL5thurmb
YxIj9GDTuLq2/gdj9g2Q/ub8JjvyvfH48x0NoPQrXfGUnLP/zHlfBhzCVxk2RZ2XrPh9WUqu62ss
BTNOxvL9lfPd/egWJBEfYp3t6Z4clWTjVmgxJzsMPhvHFUPQZeuZagHD+43QcjmdNUgBoN/e9dT3
ZgsjCe4EwJsR/bxC6KnFfwK5Rk9bra1UJm6U4R8w918jV+sNO6hlhZEChCyiSdeYT7iK+lh2zQ9p
hUkQ/WjqTWzqj6NbZehfMdzSGzrXnrDSGydv5EboIAnkE4VqfubrS4hONGaev6ualqclhFctxRuD
7RC/C1NYo4kOnPoOb52v0ERhfhnhTqKW3GtTZawxeg6v6PSQ+l0f1bC2HnnAepUhy3B13iLYv4f9
qMRBPFb0sDnXJNgEadkzcIhBJnDKJyM+4YB1bxEGsV7q+m4IBPKJzzsxf6kgoNkrpZKTJmITG3CF
61ylrQ+0VrDvNg4fChjWDeAbfbIKxAtOfwncwWJH8gHkOb58+O1i+k4zwCNKnllZ2Jzg8/kbP0B7
nqll5/oQTuxFqYVGVVK+zOWLb/Nt18E1f6Xjz964/mGeodoJc7vYGAO4HoC6kmGcqdIvCUG5ibE5
RPZsECCn02kkAm5/XR0x3E3t2ZHimDjgd+tF8/yKu3hPhQtSigQxrbAYBuXACR6WUnvK1kAPWzNo
S39ppUe2J54shS2EXqP13a0GYKuRa6J52rDykgVfU+Tom+curvVyzIU2rtxZ2nYsjqdHg0OfSNLJ
6XY+QP9n3W0qHuTBwRF5tZS8QbC28S3G26dJu0jFOafPF0QRyP1hQtZS/4Knx+9IstXrZSClEJzG
gNwRUsFanS3qgshZc7NsrYiuQ9lA6xl0Ts0EtunqZTGXzV0Qau1S1cHVTcYTYTYmwsnGOhNwsReY
71OcCDUrqemXjjogcQ0Yq35GT4wRgwsQCdR16KS7zdBe2KkaGCTNfZ5DPs8hVQwsjwf3TAI2xCgh
d/MsqidKNmugTHAEi/D/x+/JDANhSTNO2xBRXvjsz/pwCMGt29GYlkMcFGv40WQAuyU9Ps71f8Lx
4quMKWVfKyTF3kM6q7jamImYfohCwEtvimuRe5GlWVf0BOlb+SKaU5tI3bY1iWBqXCYBic1ZjYw5
HbTehR6r4nN/Eme1JkNTW48WyEDXEUWBF4sfu7ilyY9HsNaouWmgXgHk18LsYoi6DktgMPcDjAZW
BZDFqVIMJ5F/0L0h0Gf81Q0Yy7hP+SPbb0oAQhc5gJOT6eWNg5et9iZzxeqXNsK+gwOEuQH+MrZe
TvcO76/OJXed+2uPbnb5ljF52mZXoQyn8WklUfaUlmp2sbn+EQqfSPqmfiWDzwb4IgSR+zrnenWq
Q4ZQvvAKtayiq2X9txbbimJutttXlpp8SOyzpJrirjWoJESIzL7rJYXC089OEosGcE+s3HohLWy2
IybrmZiicEhCNm4EeGZAUhQ63JO4hfLVHsk91fh3EHFMefyQ5C25NBPs0ffev8ijay+cUsT0hkWr
azbMduNlUykNrXQVJmrTRj8JdJ1UNdq7rEy20psUBaNRBbJp2qDx9yldX7Vsu9izRVb+z+6AC/XF
OdcQ1ozadGgTok+/7GLcSPLQmXakFm6awshPizV6YkdUFkIlEl5gJ8Yb8fW9E7BL05MIILZHXicE
pcUDMpO1/DxnM8F/ZAMpNnMUfNisSrCBbp0SqM9t0VX1KtkAoX5WjPLcSZ2fz7V9sqij0IGK7UVB
UQDb/8osrantqg4Y4XuE/RCvhRpdq5k0eNveJAIvJLUSeLcVtA7YKma/G9quyPnvwzffgMHV/gwY
IBc2HdxkQSOuN7J38Ihbg7XGtZuM4ALcL22htHl/MosvwgsO1rN8t1tOW3ZpGy/X720qNAPT+BOi
tR3YgvkFZmQjPnpe2G/+pGCJpIrK3mwLRW9tUErJ4tQIBIAz4MdjTDjaIKWyCxDdykQYNtzvU4AF
Y6D0nPRYInh6ifbvhmF973dPqYYsnHIJtkcGf0PrNW2JGPrADHNDAPhvWT282C2sVObW245u+9k8
H8D3ykYqNFystrNvPDPzRtQcBv7Sw1w+JhfX3EWXaLVLEzc3eLBb8Sv0SItWmHi6U7JrgpBlgbuN
ug8Uab1ZbHujgDMVSb0wlN+usEdaUSmxDZx0GwtuPitwfGfX90zBXd3gmHUZzYafUjW2Kflge/sp
CIeLJ+EOYpmCF6+ro/q0olMX9SreSgVxv6Tgfm9VUlfpYOgUgA+SrFFJ3KV8pFZ3tseuqoZP0OlR
uzmjQe88IK2UxA45xDL3tyX1gxOQG+pnIW0jb5mjP4+x9Qco9Q58sgbl9c3TnSx5IVdIz5m2bTPc
e/+9HyW8GsLpKomaQTVwGIdfIpR85q17pLEOP24jid2u9g9fldzYv8GPPtYR1KE+xtM7WBH6nbZq
50BbZK76JGXUIgNSfsY2SIfDuAquJ8aqExRrgUIa+Z5B5/yoo0v00xULh7Y/1DGsEUNFdU2Wi4k4
BoErucKqit3/JZ5jh0Ia/1S3lczjlzuKV/8kXnRNFPubqMlzGumFJ/TfRpSfEK5V5o0QjD1zNgPj
g0DpaqXLL+rWau4KzOIRfW73eOgMCOHo/4HUNqIAe8b2UgNuFOaX92/zDcbNLyve124wiKyqDooD
192sgvl7+mzLfJ4Rd72ogzb5Fopc/t10muSRrC4H4Ey/B+fU7BlZvODh0BOCQbmbFbAAH4cqSkig
K3l8yIVPfRFaRhE3zNghzkehnZqPJFzUy3mRefMNyJ00v0iGORw/C42ZBOCffCfybqOZCgjW4Ndz
Ys2FsYGrOOnZABdyTsSvV2bLtCPZMTMy+DDjBnZOubKJ+ZwHPrbe0U5coXbFYpr/UIipvO7Mzdtr
eK+jKaz8dyt+KY8lh2ddC5X59Or2itJADYMXSRHAFAXW0b/Cj4H+oPmGrPeB5A3m5P2461A0Ejdq
ogclgyQoROScFEimQb1uAqHrIlkAjxpy03aOjjGJ6jqQGQJJT5wGvYSN59CUHP6JMdPsV3d2/mA9
xu9IzEe3qPV76GnOEZU6BPbhLGcDgDx70Txbm81gSlJa1ScA2hgWG/PJ+ceHPPHsiai6TwKsyEfW
E7v55pMtyZqImqZUU6sEoWzfjV6Gal7Yrop6ZoZeYV3twtjUwpDMWthot+i3iW2leb44gWDhSHY1
O6LuOw05o0C4ihMyzJA0P+dR6SVV2BLSH8qJceMGYBF1WMvK0er17f4AxAEt/twwhrapamrDo+CG
k+ZUg6/1tj0wF6FP6hLy7yl1UarIQNyRtqWrIMAMLh2uZtk9diWavyV5LAMzdECvhoaCe14uhCIT
KvqQIQ4eAAfPKGyTwpGnMFXPrHyWs3p4oA0ZuGx0e9RlFBv3G4FfgdTOnp4Amfpgdp0CMTHxxk+/
8NqmJbuWlGllP/VhFuYPCctlnug4xzGWxMc+2Qdhyz1MA7hdebibi2QfETlEi6PPkrBayR5p0EJF
+ffdyvv+5Eruy7ere5j0hn05AwjhGwDHFdzDAtKu1SOtiumYbs2sWf9dCMyVkxZNhBqFWyK1EQdT
ak4agDVG/4MjrrVNNNh6tz9nQYET9PcogRKNPka5SQgNWv1oEr/mzxNXwKVNpqyIhCKqFI/NgE9l
m0SzLluL+4qvyfm4EgCeidrqjEStvu7HOl4r+xKUx53Rgg/Sqn37QqPLgXhJl0axUCQyRkvOY2bb
Owrd04iHQrccoapER+U+lvQUm1HKG8Lx+jNk3fgOaNfDKGj+whpfTHqLY+Qe6+2H1vqJYXcLEdo3
qexeheOTKjqQSY8sw74QAsF38GRH9LfgVMF6Xt0lvgippfccj1JQxfJmus1yaNjKhCbRCSKPVq/E
zYZGOYyLTBrRv0Bp5AwqMjnWIMrlTy4r58Esq2ncTGKvg20CXHVGKg9qMyMmBwnGJBaBcC4JkAVH
Hl3UkaqmCfdect7lmItn9AGAAEE2GjL+my9QKpEtKfGPEjxzRKuaN5uEJ7jRM6EgRTh05sEF7wAK
w7Tp5uNsDmo2gGCaWrUAUnSjhiw2Z6p9PWN1Se2xVOosARMBePNfJQxoaZYOGTJiE2qn9YUmW+XT
OPWD8H8xaNtrvM6jfWIRsliYdEygq5iWd2JOGsDNS25o2zpyRamrMng8Q0stfmvOQAyeiURwJGmb
AmkOA3S5Q8RdW3VUoQ+3pG80h8reV1LHYwxsiUTCQ5c1VxuvRUixMjdyUjojnA3PIkLrhBJAFLJ3
rTaoMDC57wUn9uNVua799Sb5hb26XmGchUnHqRLoq1eKXTSaQ489isgL0TTc2/ZeP66I4169OqYm
GBXJ0IpdrTZln7c4WJYzqV7LppwKmRPRMFzqGX7q3qbUdalURqY4FJQTzWFBBmFQYO2n8TH0swaq
/bJVF9H+l0DlITMULCoL7Dgu8OxjOVIMbxMYRGAh+JxKR9LrS7vrMIDN36Q8+cmdWplZAX1KxlVM
8qGqQWZVYMFg3kXcQLgXg85PcxgyZoV/TTFeHCxAi0M68hue2NyzZ6dxeIAkHGt/Hv+mCkrh9VmJ
2eJSUA5pUAkbP8pGOFiN8PRO4ZeQ+uQyt5ivJoBgttUZrMBkqPnKdazZ/eb6imxvrGK/FfZGYWMl
6ViAWLFZPoVfTrKu7YgteiXUQvR1gkKJAcp5F7uoFoXWC8sAqEJ7oAxGGhzOYkmXb/Wu3o5bBhJS
ZKYNFl28vHX7YXyJlxNVwF0UspMCXRQ23hKpbn66YFwjXcVRV8hbDA6hBwOBPp+zP+L5wdbyLqAo
nS7rajjU9KMYesAxD06S+583RUSam54kqHdUEOoggYk0/Jx53laAnnXyiyxnlYJjInxku5ROcaUE
NVcgiLiJ098j2/YkbLSDNi83Kj2HriiOhgERGfk+7ww7gY5R4xr46aPyT9F1TKmh/87ji/a78LRf
5I5RMXBbEv1XCHIEO0/iuUHvdhVs3hKWHYr7PIXe3hgV2rLNeoF5ige1+NTqzAjtsNmduv2sy+u5
ivTJ+vxzeAdQeIijq/4LNfADvkU4Vu577lokmT6ejLVVlZ/AG4RAnocJk33+LNn/BDGMtkJjHUsC
ELQOnkXU8Cab9bBZtkK4mkmy02hZw6wajwy+4tjcrNP47cFOUeyZnRhkxnWCmBz5NO+z/V18RW0C
akj50pv9suDjQ6unrpKiUTSEpFHnVmSw97wptABpGQeDOn06fLPULj1cR9Gv+g8Hswhlo6HL805n
1Sk1pfrBTDZSZcRcrf/DGj4ScwPeOy2753MI1fC7Wn+zUWRunxbf6ELB5GH278ULoOYjdH+4f/Bj
Qbi5oLMM+brCiyKvGpUTNp4cehwH0zBWVmcCzjun784hpGVMzLECXaUWxlmXl/YCSQG8nHfszEO3
aQAZ9Nnqx5kky2q1hFgtNr1IbhPsB54c1xpveZP+PvPrBhtltNV0gMinzfwzbq6YKjSD7fBHVWCd
PSvF70Hl62PtMCI9U9PP5JvfgC010l2jECti5aV4qMDfUy2Stk7B+nZkDwCk1t8k1x2PqX0GsnWb
QAFz9oa6z9mQIcGwlJF6gJ6K9lSwXoABTYn7ilViKgoPEXwlIjIrATmHje8NBQU6FDHXaht4qder
ZyrDcwH9w+v2DbqCIIH0egiPookmGpYYk4Qkse694f6IwcyxDYbAghnNWDFcOu5t0OqqSWtYS3eX
tsFC8SMjlbSYzhWcA5D17lprYsY72E4QVcUcrHHfcL9YCvPgAFoh1xF8OrzbhIDkpBtOJNkwtIX7
lcAwEdRQzAwHh3JQP7uiKbCoezsFwfDnUAUWV9qpPz6OFrz/5DoShdTyJWgu2A3ruPFMn9owiiau
HfNWPoclt8hEgFE++Ya8E+JhRoSsedo0ddBJpjlwA7EtTGs13VrrZcVQxLMs9XIYwDW6Gn3hRG4z
ePdiNvgC/foInJlFUh0+dO/xpZ4mt5tYkhGVrEE/Z4G32CMXSo5GIjMZxad7IWmfFQCZ/I4tpdHB
g7hcXuSKHIMlKxa57wUthnSCSEURhAE81Kd5qK0rJyh3yhtiw9emEPjOo+zQWrgkEm4n4bUMsU/r
1yufOCEikiQMCnOHdi5qlRwTfjZ6DkobbUhOjy6UVBfJHpNoB74gcZTkuN1FPzF5Kh6k4jAGTlE+
Zt/qXhX0TPPdVqLpJk1mCPX6kJgIyoimRugMnFFNbi6uv282gLZ2Ol0MBu/Q8GVxX6LEhWO1Azq9
wzus0WDX9qP3Nevnmlk1qZakIdj1iXTd67WxComucRVR/uOrYOO5/PClB3slDqjANJoZ/yjkDbyG
A6dNepf7WAbQoV5+CyCQrrhHGHroQ0Edlt+g5nH2QWt56o7UK9HLci6PG8tyUmjJw78ExjLxFcow
l73Brqe9q7Hp6USGwjduU4M23UWdRbQaWFr4snmVTuqwekgr5ofKBmmcYpjrkP03LfpRugsAtiUf
mvG5ft/9OvnkiCONDcFAq65sqX7e7OEayY44PxFFlqDLeoRwekX+el84SSyM94yKKt9SBJHhHog4
r0HFhYhApg2ODgarZYCvCq1nopLGlKZqJ6H2yObFQupaA+eER7KVhbaS0dMfi0bYygR0J9uZtY2n
zDJBoBYC+OSyqrESD33//EsjW5174J8l3hk/KS0Av9MQ258KHF9zSW4hBQsTYbL4yy/kzOqXbuAc
+qxwCPWKp/kX4yjS+umUY24wv6NhvwTivmO1hDTYzUjcJT6dvS6UtnCxf2TEVQnJ2t/YJj3hfnR9
WboObt4Htj0eNPSJQIXrPuJ6Oal/lmLF6MjkQh3hHyVd8Gqu0vRcX9yVR8+IyCtcgSbjX1X2KSZj
l2RpokGuSQAguh0NAhhUke1DKYc1qbVGKqplJgBlisxIjkJdTsblVIvA7xokzlUHdtpOOChLW122
MKGuF6I3R217tN+lTfmHPnaAoz96AflDaswNaOj+bFV3AlM3N/KwGMz2U7kboHeUrp1snDrKf6fr
r58HQxQUEmsWGjmpTtBW15GgR/4lEL366A6x5WpfjBCUZbeq/+LvjKRLZCj8vPgBe+Wv8eLXI5SZ
ON7E/YMgCKaRnDbQROiQrAoRbSULo6XMouSY3DvM6zppv52WZYViLpWGDvbwRkU6nY9v2JjOb1/5
17B4aO+XhoUjMzlLkJFlbimcthBmHOcjy/w6HPvkDRmcDl7GVhIfs7yYJeMwueDAcTcdfCEmBcX2
8T0VKXEMrm51rQKksdDB1Ljfifyhy1NlPALJTVDFI85PsTN/Lulz1+5z57rkSqLAos77OP0TJiUu
UUhpLMrJWOyCU473naH5FGq9jbSnjk7t6ErecudS4wXYIkLHJtNpchN2nrmsGZa6rPxilNMAyM8q
mSiYFPzILuIbhWvC4ssZcw4zKnPh8PFg2USnrG1PlPpNT4BH6O0GhFZ3q+97yFjvw5qwJ32xv3UF
Z7vhuRW1YKQ/ua0HRmjU4OhqK+yO4PHKoCEc4MBfqxbmFKxc73Sq20QaiY2k4S5ZkBzzSo/w7pAf
SiSQCr+kBvDiPNzT6Qaamikqgq7ES0zXSCqcJfrlFDD+Z8X1UBPLbOYeFj2Rl2x/hnHb0+JxWDZJ
pO/VJPRhH/+XJ6h3PgX84W4hWLSmp0ZbrRgvuFdWe1PYgAqn+cqrT0Q1wAP2OIu7zMYqTV9CbYO2
S4Oh7jvr79kBz5FsyD96LvzmvvaB8EXRCdXv51mYiK/SkKuW3qVGtuGWRRNnb7k5nARP3/6CIMHM
uliD1rPY6jgijwOWeVyCS4jNCR56U6VVafLfiOXoqeUi2cq9YUQ65XP/GxApdvy1S4mXDjgRBZbe
ETe8/wCOeQF127iP/OT2Jlc2p0HRxWWYVvC6S5/BssnGDUF9VWIRYJ4SdzadM4HhVZukhFMDtjTn
zvRhbP6doxuKhGXtq0o8RXJFY7N0Cvy2LFS5sH6xSUw1h2jBzjWLDImRKd6Zf8FQr3RZbmXvNQqK
0G3CPpZvgK6JPM6CgMXfOJB5Rau+TxgtNdmEKvPZ1mVO/TVmSAn5IJdwbh+BQ5H5cXqLxxNPQDvO
+60BDbvAtJ5nAGhJftRp1+3LwVZ3hvLxRegikqXYcWxyV3II8Xsun9nQEt2eB11BPJSkWfHqbObg
j9cyZRSz59nQfEktA5c5SBSwUn/rhErj1m2Ds2LT/6iw+Jm/wwwCZKOQ6FxUC/jhhweJiYeIipS6
zHeCVtvxIrLVI+ruuKmU2Ffhlv27hpRj9dBmb/eqc425Y9yHQXllFrr+k92BAlnuD/CCDYp7UJbU
4QSGOslD9VeCT4wkTO7FdSQ8az7Wg84qnxz/LYEmSm3bfxhVfqyP+IYTzDiM/d2JE+qrrsxsYDQQ
aNH4BcnoMuqkN69jVcZZlUP990g7236D36hMh7GNX4+thy5TgsAzNs6Z3772Up8OiV5eimkqljsN
EbOkT+5ml9ONs16lBoYnSZqPrl5TlhqBqm22RNU6Dk55Ir4tuurgeqjkhG5KOfnEEJSl7ER/HFlO
Ga6g20nV27Nm16V4HShIm3k5C1v+j7L3/U5CVsQZ6Hz3xlV9Jjzj/lLQBMhXbpfbclDh1YPe6j9C
+LaJYpen5/vjvn0MoLOZSAS9KoXmGIi6UBG/VAkJNrLTSY1IvVSuBQWGB5NqOUx9lCMTbIKBJBNT
Yihz6LxjlH4Gbk/1uqPGCepMm93lq2k/Qg/o4lC7iR9up9ZALNGvvqwQsRhzOja42MKiMmh0iTas
CIHImJZgCVoC5gMa655erIQDXX8BNOgg90KoYKE3KdKaPxxvfDCdON8d7FsuAFAR2nxkWkPWWaHX
K69X6u3LJTC/IzwYfJ/bsbVC+aobdSLKGXcb4mOhXTqZjshs0dIaC7ovUZvz8yyLxTxUODWGpLr5
CtkPVEHRNNDtwLgVjeyXBHmXtQh5Zw+B9qEcm2tOOZTP8EgKxqiVRmfwYGz/bukSBy7L2ZePinu6
1c/6sXmcqbcw6W/WfGvyk5F1qZDtdLERZSMvsCm5HU5QlVlZyhOzSeODn8R3Kbk3etUXnOBeZLQp
AOOItgn0CuWR9uj6wH6nMYJwYUv7st6Hjz1dfu4JDE5Mn0oPzFtmaIo82JAtqoPQNA8FGRW21QOt
7kVrAqwvjSCz4vFyeIqSvCK8ZDU/rpE0Lpkh4NiupJU69m3Iq1J9ud9eop+TO2xRAsu1Gp/x1XS6
xD43Il4SnIqwQ+wzSu7R8BfgK+WUP7b55mwTB+vQO9rLeawsJ9qfsEftn8ZWDSkCiVGH9jM8wLBt
W+K2JggfUlq8DgBaFKqpW+Wimr3kgr0A6WjJ3su+I5g3Eq8OtvJf2Y8xsaBh/CGeylGaoiCxKUiI
pGm5T/Fkg3QD0/xEEIxDGsdCqTZR6isxKogPQp92xR5Jm95JY8nlysf4z67DCiXeVN2Kj9Rl2WNR
poMYXcMGBUTYscV8ih4I57bST7GjvW2j7pvikR7nxtisGbkJX+zu/lQEvj06pGEpRq7+qlHMcisb
+yuLKzt+oD0dfd4GG7Iw5ZsSMms+iuuVDkQznqA8MJwjTLR8qu9/5Z1egQNWt/IGK/RO6xg5aoaP
JhfHwOv6xzwZl56/D4dHjoPI4nK2JIYqyR8hzzSmMu/g/9n0BvuZp3iGJJIwnA1Gz70YOanA1eeP
f9/3Qvc32jukc93EMHNaH9i6mJ486/sdXaS/riTJXmgGACVOGKHR/o0S0CUpfXFrtaSFCWvWa7+X
o57af2ZGA7T2Y2TJDvoHpEpgzH5pFY/FALoKJzhDoWkdY7JDpfmkiCq/Db1a37Q4yoUAa1Lz0k4U
bqpUH1/6JnQa0nmdGNJHJbNSDTRB8hU/dDtNsTDbypDM0+uvbDqxVVom1fqwsBxEFstCUOaaglBT
pcogMt1r0PPn9b5+8NrigpWX9f27WKKN31Y5W5wAkUxeFpKYqZ3hJyn/kdxOy5qJAyLpVHBgn64N
2HTWRekH68iQjAUl9BclsylPD91uWg5semfNlRsOKzZ5N9N5vhLxg/U+LVE7BKU/etXqNPnAZ4YF
y/60+cYxtdqRjkUN7M1h8cVAa0idsebIudyExFjJWghvKcSB37qGRiSBsEM97y7vsNU2cp80Aqcr
Wwuv7uZXziGC7QCumH0LXCys3mh5pHPCWJY+kpXx2iY0BTeW71Mbs+SeDlUqtvHzwtFvHL/oGecP
1sY4P7BaFlOimQukdCGrBcWfl7yF8wMJOCgewVJGOXAdyyJO/mpo30jqmLJa98ff1USicCKVPhBK
KXfl2SpLvPMVhH0St9K80T2IDMfkjMdMMtaotugze6GKMbJ1RYQZvu5HhqcXiOAyaU5w5b8NQwRF
t+iN7w07P4XT37OJwk8z3dbA/cKOI9FuLXbUkMlMepFkiOl6rKkycKPaPac7NIA9LqF0OD2RTz4y
1uYK+IToNue0jEbZ0WzOjyFqMq5GplUqWQZTpmsF5w3z+C6Q4rM301pJAew34Lfwy1G+PjM8Z+YZ
PPEh/SLlxK7b/cqxqbdhreUBTv9NNzQXlmg7vOB/FgYyTooP3yYNZsXsYtWdAqrwwxCMp22Bg3zD
u9KBL5VLhbAS+RidTcpKfgLQCsasmVewQTTjIFK0G65tN0d47mHFTYNNx91fdyADbWbvuhCV0vJA
vkAm47EXjB5DQdj0eowDUYDM3fL8zwzvIOIVQFkNet2p7mJcbKNz/nMRxqEcKoXFuW8FwEKn+eix
r1r71K1O1fsF5TZ5N7D64mVfk6bRr2DlDlhaNljpKA9+a6nmuBiQctZtibTEe6EswTVAfR6gySPT
+KLoxYWs1nBM8qnR30BSPFa9rhQ+fEqh8gYLcW9hjBISAdjQebYW22pI/PqS4PJP5jvigShTJDE/
QE3I5eatb4nrDBoRDRYHjTLHJAvfJbOw/oEeMKPwbctEd9045F5xrUgtLDP9MlOPdJHh9tB7u6sX
RlivjExOBYUdPKoSqnACLhrGnhaXRoSQ+4bfoKPY1aaxW5dTNvC28QDP9G16I36TVJ10o4tVOUBA
YaCc2m9SvOvPWQnVBQULbUgFRz/81Idwt5Y/pdp7iSGUg8Ie5I0prmwi+wQu/JIWdqyzsy8dfIeM
fZSdpALjTMd57WIErzwoURngmcIg2sA/sLe2tECiAP+HvJYA5i9vKUErqzU5+gIwig+IqTVTOu/V
7aP4tmRuhj6JkfyTIhAq6Fy6qsfjByctooxbj0df85dLa4NhOznU3ZmTNxArxi/WD/Xcyuo4OicM
TjuKvJVykmHFvB1Zwmjiy3q3RGfUattUN3Nbk1n+Yi7C4z9Z/wMi2g0SGskoAXSFIpN/ksYe9q0o
ZWUZQvY6xvE31Y3X26ta7fNDEtJRjcRzlyBe9yrF+/ctEvAi+RBYJJ4SD533xRFx04zhEtSOqwI4
nRRY08w9yKjnwsoL4CgV2kbfHOrkQXJxMYX/P+GFXd0R1tqZKA9Lc1F4r/uvIdgv/PRIaK2/cDAJ
rGF710LyIMil4PEmlDD0tQXdnkKd3vkhZIOdYESg5eVli0pCEQUEVYgeFTxZB7vp3pdqyCTLmrg/
dm7lROMlA+nqH41ov0Uopp6j0D8etuamWhwzVqwoOT7/xJT0WyPxgNK1cn727lkCOg2G73HR5w5x
oB+nwCk/wZ+Ke7j9R3ytGo1olXOjVp8uu2zqIpYfGsIbvW2ulGYYbQiEm482hWoZQcdobGWsD5hi
YkHjgsxYcVGUMIYKcPX31JZGZZOtFgG1/uqemPYwTL2D12a0FDyUFmLMMwgx/xC6GH817xbjte5/
I5mYARwTMj2r2IV7hrwMoAOM1psWFm6dn54ZvAH9SznyRJVg6BQfFBk5DgitOv9VOcmEP5pxijkq
rNrEpNeZZjMQYTGgeXNGWBAVrSkcge3VTY6VChIFwhAR2FeOITrRLgnOCtHt7LMFVKSK+ffsEFUx
OX8ovRza4Ej8xEL1rHVV+w0nE7x+zIonbv4dih+T2eLzPd9oUogjfLgiLZBxl5Xn8gCepwl0y5cz
Sxr0QGqw1qLooipK2Aav0kYyDe4bKdqmFMZ4keRAbphoPFALn6RKaW/TNuSZrGoIHQSWV7pqaHrh
EfEgMPtfrBuypeWq0lKmaVOG/tUFbj3QQ9LpaFxtveQZf58pNye2iX44Jn4+v6XXhDVYdOl3CuFI
qye20Rfdy1jrMMfh6f+utTYR5Q531s7c4b3E5Ni4Bq1pkIwROPyhXEVncrqkrtQcK/Tz2SH8DECZ
3QqjZhWwsFsSYMu8iqOJ+xbBFQOhmtcHq0FclPAHIcn/GU1UpIeZctxD335Xu14uhJVElJQyiued
Y0serkhune/XTAAdwhU7VXN05qA8tVWWbuf4xmPGlt+TajA9yMAo01adk8KLIH9J047SWCERBUT/
7IPOLzOPpM/5Cz1E5gc7SVjjT12UKmHAry4EFu1fy4T4lryxv2694Qbm5oH/nMOgUMbEzsRnUfQd
mZzd1JjJ1zRPKL/b6ScuYb2t+UDAjfLOXQ5L4R/YgH6i33ew3SAi9Py1ztGpBofmBGH10u1bPd+c
nPDthjmDxKiT+h8SKo0wSkz/d63wlmAkKvb0VDm3HwdapMM9Zfdpp6TB12Kq0w3p0TIFRvxTzNWr
mURDmhAaQnVrt4QpWFPoo0I4CTIT2NdR9tF9dHu1iaz2dAYhFtZnE1TakxRCkGVtaLGgA9ndsJGd
KJ6RtGngvOOiYDuWFtGQ67i+nOY8tfy+V+kofgZJymBdQ7Lx9YDX5s9rAHfDdas6PmPqOfM4ZkLX
+pErw0lMHTmSGCO8DZqWba/RwU5wgbevRyErVB3qq5l2qoKi+RdRgAQf3VPYmey5ZbZzdODNDujf
Od2o/0xp501ikJZ6zLxGyLlAS/230UJjSSF6MU1h5xNKI+90iK+jqdnyd8r7dfVuWv9QNr13xqng
0a/QPwpE9u1K6LLMChlwSGoVEm1VDXwy7ePXICy2sDVI24AX5xT3Z7Q8QKTbGfADvO/U3c0E0h5p
kMY3CzRjiafeRROyM+RgEgDBxhk4MSFhHtM7HZkGulQLZWccKZMO2dgRJnpfIVhdSlCX/aUB8/oO
u46dIpyRxTgeRkGc4fSiOOd9FiLvHOoSwMBYPXzzGFhHf6Iy07tqtrmww4flSpG6tU6pG1ZITuYO
AAnsO/2VEDqwHuTIsFovs4AnLoAZps55nOYCWqsdCdY9PfAXhhjfNoS3QzD+idJQgxkseZquep3I
BD3HAnn02nr+pDpyI3iOoTS/6EnZHWCIPYx5csx/+M2zbWYOvEM0g7mzTVQB/3Qwe/abUd3EvkkA
kbLrBQu0BqNh6NAnkcptzSANiP4jDhj37yUTQs4IgpmMbiL/kbCgTiuxQE08wT0yDid2/YV5VaLg
3O8MDmK/ivVOkVxtVrNhk/dY/gTqRIhg4fTDL5MJRkNwtm6whjZajTfTLQ10sQD5NREazAoy5eJq
0iKvappG5DbsnGym/kQv60Y7ouoveJ1eJSQEnvRsoEBZFN1MO2LMv1knLUnYlAx52vnaPeFWw55+
G0LZxU7HWyGUVtKo3sgdmT7FxGkUlee9kdK39sq8fSxTSiPiIQIiKkWsf7vbxqYz6miYOiI2y5VG
IiTqfLNCNNq7XsQS6H7Ref128XWX+LVQ8sdzlwup8TaYFR/aCElse+GblAQ5Buw75+zfdlFaHZPQ
7STi7PSjNpBQMQtMaWeS0NmwCVpW3SQfxx+57CK4H7CP36EjAjxw6hK02r2r0NKK4oeEfjwNUEFG
ZLGiMsj3BzaLijhICFauntUqAa96CmDxgutydQWwfxfUj4a6B+Hjiux9w1fm+++Mr08lWZy4ORse
P3odL7py2k7a5pUPyDsi055Djmw/Bnta7BprcZIpVlOeL+1AGiJv6BuuAE0sB+gNM4FaOyX0OnVh
6SxSEYnMuSbhl+2J1c56KeTrWE7ZsViCp1W/bDWVLmQ4RKXOPZQAx03PZWafxfJzSo+t7odqhdtL
sNL1bnilAtUoMaW0mBe4h3DQipjUy/RMlOMSvJYd91d+HPFOPnaiT3TWmAaK+NCuGKDvtdpNPbvJ
Rmdtx+XamvBLYKHpisy74FLaGz/pOAgcVX5/VIeIxRfi/x+TgxTLjXmqbPHOk9e+1UZqZBcgMzCK
o3KR5ZyHjkjKLUZLdwx3XxKsoda/zXdtjkLob36oPdOQUlz1n1a2OSLfw5ouWrsPqI2fAyHkyxOw
TJpUxTEWmh6MlEq0moICB2K29coRi5J0N1fRiV52CGcBAkRh1x0Z2Jk5T9vWjzCBnvezdBTNpPaz
GRkkmcBl935wOd9bUjDZ2E5WExBq4rakYZHAQcymdIFYwGLP2hjdU+ep9KcadpNyPrjkECLoBx+E
Q+IT6gP+3+Hp78vu3Qk912OQ/381mpJNO8v6mVifjwA9vM0PudAMC6fmcFrwBjX3RJGik8pBrNvC
TLhObmFyvYZE0SPcpQhQmLqMSuymmCrUD30VtMr53hHhez0+ZehHdjyHjV2On8FgWSuOZKPrQ6An
RrsMT9x1TtlZuB+v6Z5Ob6K8GLrYXXptdZGEBHKSgeciFqtmi5F9R+O1xHdE7Bpy86OQ6PdDPlC/
4l5D56jjIwIUJCpahppV21HYJriSiRWamRVtdgfygZM8YWmTG3/WidD+wI5f7lMwX2g1I0RcPZP1
nwiA0v2VFgME5AsixTQeTR9SF3nnI3SQdZwcJnxW/Y0AVrkz26EaT0uzJO+BlZHDlGHpQrB53ajK
3jWnf57pB6c3TryzxuT3AkUm0dW9ej80IDbkzGT9SpTCdNfsC5xH+HxZhhaj5LsI0xucFGL0C/dJ
8NlIIfSgXLBryveU8wXtFPqw3wc1AtuiQgLpRIt1dOuGCR6hVmXV4WpKfT7mDIFqR62yuo+Dsw3j
pIC3U+6+BuIt52/4yuiZYE2KO6R6mB6VlaHtOatsOSwuHjTFsBZONI6oXeEDEcUCmZOA4ho9OIsC
aE719jXMc189gaPoXdlc0Vh4vCk1OaoHDk2ld+atNdBMoNXS71bFpUOhAjBvanmNQa55auUA/aIM
XU4aJEch/HFh0DKk2icdAuSoXXasXIX1zgNirgftOTCoU70un9LjN58ihpkP4XhNhPsAtcK9MNwo
UdFXQBFSZQ+N6zXk5foHYkSFT97l9N74ejMlK8MS4wHmXSXzXXV0K2sdI0gTrFodunVyv8Ol4c8K
SK0lY4xo9ZvOexn6FrJA4n7Lr78PcaYrvMiRCP11tLa+EPbeqvFeXQWS4+TOj4BTMTO8VwRwc3us
+ePlwwtPBOrollTcEgflpc4E+geCQZ1NP/8BNnb2Zhc0khay6bR9CKn4TGxYD6H8fJ9+GzicFxX6
WKAVbW+K8VwBHFctuHBuO+9guPHcLh+ro2M7ob09WSlVCZnUTKeHw2EnnUpZkUddlsewWwJpCd8Z
4wkcIiSkpWJKRb1nYAampeaCuFW/1l9plF3MPZTMNEHaZ/uE+XHrCokCP0dDzK/5crXfBqZHzEtO
JM7efOhRUmnQLpOjS5E3HAO8tenibvsb7L2wH61Z49BPLlgD6y6lr6uW8TaPBNxFBQD6vMLxHbi+
pHWiXtk76yndJT49HCcRHTWQ7+Pm9zmPetcvgI2ZrFihkYbTm3ZXmODM3WajGjfLTOOacBR6V3kS
t/fHtb/d47gQBiqPZtuq/K5QcMGN0DjibZaXjH2NuUjkmbUvhGgJhUpHV51eqsIQHdlc0QPTecxF
jpExQmguTkMJfKjxT1DaOdx6jGnGit1mE5X2PZpd8ZeHz88fa6AG6fD2AKcfmbg4l7/6m3oo9sTG
CYEjpm1lgc+VeMFY/4h6ym5kTsmJr6BXugrSSh2tnsT6A7IIKENoUIdXfjkSjkikDs8Dgv2TOMN7
Zps0/W+fNvtS8qGXtqbtONIHqML8O3NkbslRBCR/KE9jSVCGd1HNh8Csjt1k7Mlc4XMkSoVRJkuO
6uuNxJBmZceQdaw9AfqyZX+Zs1R4vYSM4940Fx8uOaZabcYij37JK1KsFrP9jH5fbUKOfvYqs5AR
oQM/dBypoDQz+DWYGzzc4IHu8gTlInWqofK/XoJubjpMIWvhzhHCqB1bKDICLhL4F+zPgsxjJ1YX
NdyKlnBlx6IVetJynii0ecLjKMS7dABaaG6+nYk4xkNKEy3xV+yX3jQWa7WGV87VC6J/X2vSB7Ig
vTZ3bhTuUlfy+sTIv0adAyiYVRrprYvyQaAql+9JYblxdAnftNF5Bqifzuw0zHChxvH1d8wVjoHD
GHwSMLKKE+90UgAanZGVp18/I91UCGww/08XTMs0RuKS85lBDbuAuysJpE5yZ/lutvF2fWRb+bz3
e5tQ6OFosdW3ufQJLPDpPLC0U3qtyZ4WUKL6GAhdR+/Y/3LlajDJzx5I2EPFqbIDCqTi3jhu6Usb
hWSW+mQDyIKKPz9l1eZApo+Ug6ORfyvtMPHyV6Jmbb9l+OhN5SyDkBccIgCsB6YpAqo6e7zO0it3
+TuFeqojzhb7BL68FnRL3WRHzUTQqJ6Zu+ek5nrVZ/vua12aenR7sjig++K670T0F8Vp2xm4cJbk
0ym4AgG1R5CQKbXJAB6G7OhdxIGhdCCsq0wbbVgHaXMBztBg2hYRQCk+4RE10rj2wqNi+DHGktB/
d/MhS65zw9ZjagBnlrWxDn+AF61fISd1Ztp9fgJd8JJfefWD9UIcsxBDavzpwJoVFuc754k7GUxV
IMa32AWzmUAPXdya2G6E1jF4GmFQnWGBa/E0j7QwF5KsT6zHdVzB/r5m1HvYuCipx6rYiwi7l9XN
yCprNs2ZMgpLI7Qm9idSwAAyqhKiyLMsZwA/I30jJCOQ/8b6GxzoNMitKWkgIhBpTsp4f8rOz8KJ
q/HngLIpnYN+lfpN3valHztnW5HxutJjBIvJr0oS4KeghV9RZaCMwoFILN6m+fFsDzvSKVFgye4m
SuAaqUw0H/9ft6fzOyo5EqlNYMll0YL6N3vRuIAgiDGrdZd5AExXRvkd+Aa0qizr3sOW2naAhzTq
V2qbdidnW1gwTfYXG7fCbNSn2APQbEpEBNzSF+oMuT5KtOxz+eVW2fIsNURP66VdtfQDgjbFEz8Z
1WrRLLFY7KFlJy5BLJUymzlaZJYTvIVmSoqGmiKOnO2fGYfjyVJYtrDaYla8ADH1WmlmHVao3SPI
qLPzWsLuXmWOHAh4GV+yJOJ0nprIDDvCpRntvzIMWceyzw4Ddo5nae1Gjfv+3CUcdrwkgktub17b
52l8tMaY2H6L71QJUE/Msei4FxWGBZwAbSZAWcuyKXPZQOExz4VM/kaf1/HxKhu60FZgfjLkDF3O
FB/wvHC3YyDOKTM2ZDkaJYWEA4Pz1QPqLylwJpC7RKzuOfNM4My7GNeDP+oZw4sjpzTi1INy5Dui
t6oUJ+rAhWhj2RZ3dLoKewrYElUbIYK+mS6E+MIFT7dh5KoHJ9K+iMN6VkcXCztOz6dCPQN2VT5G
eh1166L03sGRWmJbX3o7rIak/vENduvLeVDfSvA5rzz8Z2PquKXSypnzI5DuWCO7THy66sVw8Oq9
WjEk50anujptfa+Wh0HgEVylo9tTDVXCLyEcv5jUOn+IrhNwO0UY7CIr0/aR+CBWg/5K17/o9ufM
7Hm4Sjr1xyWaOvLwRHI4rLNprhrgc8e1MrO4KV5tfNNTqhMxSKzZSOp3nE95op9IwZo/nJlANgjP
GqV7U+AR+iagLyFoEpczHRf8BKdW2RqA9GD1kCCCxTU5T2HCqYsHLaNQ4S/X2Bhk7ebLaw8rSv0C
OB7hOuC/RzSNiP+0eoRxsfRgAL+8EUNlCR4W1aZo7qrKsBYqtOxcM2VLcNr220OzIRUhKyO7uGMX
IuJfDCjy5NVixfY0Gq9ZSBRy7HyUSyEyn8HJFm/q9XJWVRkb9vIao1lDCgWxHV2W0gzI3dMiN/Wb
nnbE4srIpWtDMJXDLLp2ZWnI/zONpoHKM9nG/Q85TQKp70eEvZq3x46zGWjVuQsg3Qfw13Of+GVw
T/PKS8Z4K4PWX/covAp01A3kjquwyrStNQFPeI1qzp9EdFtNIMqaz+NMo/6zjfW/Pp/A6LeVKNMf
U884grfPz9/vmbIXlPo4Ab/It7wS9JJVS0+tXaInESsFSlIosBr4D2XUpcJ+eQz7PqokdeS/W+ra
z07tar+akzOTey1ePpwCyRPhtl5KSXQvhnvxdfq34GHryC6KcOh/mw03PkFSdGHEMvwnNg+LBdMu
FGKTfjw9ay/hVGEIcbMV69eJZtTfZh8f09/uFeog5a1tKf2mGNyTSdoAtrUYuiVF2a/8GBHHe2yh
Ow1QQ02VE5fm34aO/+5jgD1sk0AKNLOb3otnUKPFiZHS27L/CIWTKP/HxgK7pe5BwmZ0yxu5/DRw
tbMxs3N7Bvo86HUGtSrcpuQlIAmRL8gLC+x7qE5wIfjJAo36CbHCBpV54gTx56o0s8M0M39eitXv
P7Gr76EFivggI1vqD36Hg9ldj3Uv5sfjEsXbc1JUuusTH9caTTEsQRe/oEMDaWtZgst3F1/7u27E
iIZAC8NJVjShzPUujMfA5chl5eyjoFpuT10hf4PS5m0xw06NF4Dh9V5cxgkthMf2b8tVMGbI/YF7
h433/DrMqms9izSUhHPo+lW2O04SDRSoSy89gt7A9BS7CQmsaXXtO6w/N36xoWUYfbKnZgj9anP9
2MCJdWneZaDenfrNnqWA5BpkoWxmaGRo/2d9IzBKxdcDQwyO+EhvjOgpkNPWyBMTjBuVsi7B4z8F
bfyImeF4KwTBu9l+CwMKDVgs0zHSeRZkrXIJ+71yKhk0TiDwaAgpcMLMKzHDPmzQS5lUa0C6DJYy
BpH52VH0ceOw1Oq6c/aJ3cQsIms1sfpPH7YSX+/tFM0bm79QiyA+qKz4DsD3wK1lfFyzAQGuvkZI
MuCZG9jXrA/pdmnR7Ynf/57h0QdGD3Hl7Ps6ybt6vGXeGVtpHPF2dcJ7JdSoDYIsmXPK9+YKjuKS
QVoHW6CdH0YXXiSj9lBxbrKpllJV0XSaRVPLJ9Jik57qifDaXHQkiCJuBpeat2Scnn7gU9bs5scU
nCP7X26sC9fA/PHzH6kNkliEOU74B1dhQpzj1ePfKeLFZr8vo9wjp6lLLLBKeEpqp1vBsnG+fjS9
ZExNoQqWt9Nb0jJ1tFXDKFcAdjK6WgwVEdIxQIOM1O6FVjF1tjRQuQJ7HNkxpBt1l2WsjFLqBSWI
vbOJpO4sMjAY5zSLWMctQL27vlr0nkkBrNXOZlipmpIrAAsRY5z9o4G7uVdUKP5McX0UEBHMnRXn
qMh17J4Ij7X9N5kZ8Tbqgmvn4LD89kPfwLxY1Qt7ifT02OOhQPZ9pJxSVjzAl4EAjynQO/0DmSST
L5tMH5pFL/jXXPdVwcZqp1OCv84ff7TMd16OCttb3F926eDv3eb4vOAlBve1ru2yGHh1pW17+zhb
d0XCif5r32gPEYMs8VyPP7ZzdAAM1EYqe8e1NiwOgTe0oYfWBUPwQIgAOiHMIcmM9VM2k1fee6RW
ICjIvIR8yN2dNIIFoz+MfEB7Rp60ErMiMTJpKcgeFnMJl1tHc0hYekFGFAyERmUsFyGfwDN/L2ih
7bWMMVwldj97UEINZkflfZWC+9vErmFKTTNl0ISBiiGTjGEntdHJm1hOLofNLt5FPbawqjqgMLEX
P9gAJiqDFgfu1csd+44jgCBY9PHVYOLObAQ8GYGJvCchCr0dL3gZ1kNpn8OY4aHm5D66cQKSpG6N
1wzGrLmXDqsOMbrBI/s9+Y8+ku6A1H9nsHBmDL2RL9ObsrKhIJjY9yNLkc1Gt9hBVedx2T8YtatL
7LXdkX2nmfHrQrcaUF978TxzBH6JBtuSz8ZIPCNk3JWGJMpa4vm4tTDpotgoIaZfYdTdDhFpVlAx
8xV3XCMglJkOXDVbo+dGRLxhHKWfcB3lOjzCpFLx+St1Q4m8XO+Uazn4xODIFvwZtgC3H2/AiPej
Xc6wBwWeGRKqtwbW18XvZ0REliBEfdihz7bTSvO7U2JXq5ZXhT6Pr/V9PN8OGPjEFFirJDZpBLj8
AaNwmkf073dGhaWtPPeEpFQexl/EUmGt0ScELKI2o5mD93AHxoBanxhIfgRdxFLu7jUIUfNwtbbO
awRcs4CcTrxCyvz9KI5x0nGpewTHWZinRMBD4pScQ10PSvi/e7bgD4PU/Uk+AFwrqAjBLlBxnKdI
y3bmJ8i/TFyvlxzLc/jv68GOMV1zGr2mdsO9ypHKGxHfUSiCm3NZnjHXl0PVyxuNoC9I6PbHyQyt
+i0JX8kQ4f9diD+bCVcO0LUfrSYVi1AgCZzm7yoEveYuTR0/Zy77+h7sZLUJCvV9CzOad9t48suz
nrdPE4DutZYCCVZQuAqi4v3sQQIG67lvb161S+hrM3/1LdQbM3aVap7ywtJgHY9YmpiVydaM2yLE
vXy/gjwBmfuulVMxreUQKgdMuiien1We/IIRNkQe7BBHK09Y64qbgKMjbzlgDx53JeLETG5dmTnh
5SpRHZQN9HR5ZoCOG5icNQce//12MgW2g92CMqn2uCK8mYUf5y13xT1SbIrfK8rLp+rVDLS4IkSq
ib5EhuGvpsSVIEz0XLYvfjPPmrfCSv1WsdOnrPwImWSFp2KOTdjc2nJACxZ0nokTVghSZCUWIfSG
jGrYEnyyyZVAK6yMJakg4ZFv7GeMGI87buFlYWK/ys0VuhZC/BeAlLz38LyZrAtJw65USnQORv8Y
+RP/k/ZK7ZwnTswcg12VasHv+Apmz5HwnhkKfBXkKjZcM58vWNxZ0tJps0kvVkh16jeGavYIz58W
J3BL6LC8FL0BY2mQSn8PwXmmfXSRhOvuordk/WKvXBJYtKQrvilvhUaoCzDWckbkpFJKx7N1yxs5
hYFFZpUYFwKbqvhdvgn/2N7kr5DzCHmMHMHmgMyM4pGBRgWUU0MgBL2qBdHIb1IbFJeN0WcfejXc
Jm/UI9NZzxH2qeKeK6+ncINihT8UI7kThDx7zobxsvlXCxZ2Jh3aYwcNnD4wJt534p3LMzkjMO5N
4XtLT+GZgSD7mppgrJh1QRF/ERQs6gWnMRa0v72XTKo/I06om1yE0nPHuxda8Y5T138OMkRRSZvV
Jrc5s9H5OkoMoSxB9cA8Px+jnlXp0j6FbBAP16dm03Z0bSr/3jYZvOqvhPrBTJr9plra2Ugxgp8R
6fULaKaD+3hZ2mneb4fDkdlqaaRDH/J/oT25w3Qw254TmFiOrnei15kVLuh1uD847ZFH3l1b6/zS
7MQS++6NDEYWUkPc4gvvxpBRn2fCVV64SyJHKGjcPSer8eImvw4ZX8USlhYoEQIIwiYg+jGJelh0
kdgSiFSe2C0J3ClJBJhl9VU5xq5qxed8oTESSGoFDhJwkX5KcjGWZiOuIH1ZQmO+fRRseU1bVWIv
6S0sH2UQL6GfRXfRg3Rti9qcYTtNZGPArMQIgTZP4e3miMyRp4Vz91qb2klk+vYJoAMHhGOWC7Fv
lj/Vpx84VVHVXv5Xzw90mUyYmFYbPu0HRscPk7czuCgPPrLAiWHqb7hLoFQ3OXHnjEkjrYjaL97K
/xG8RDIQozrHcVkUi1wiaathgnZICl8VPEyS8MVv+pFl43rCOuQMG8DJe3x8o7bznh6UxLZjvBTI
B9juze9HXvLr8ChyfErR12AGojmI0JNnDDG8nXna80xY0XogDRHX1pStIEJ+CjWlWj6088bQVRre
5ibAaZuJrOPfvHK63Jqyw+xw1Epu0KcCM/FA7XfjNEHADEoPpwOhvXPU6tEYT24VlWJaBwIJDaFm
X5dvRTgdHTl0uQldhzpJ/pdca7ygjX7QMFjJCIK4v7XbG/i12iRslpklqSOtUcpt5PU/+Xk6wDPO
+Hp2wKn1I+NCrvSobb680T0YGY81rjtl/45rmgyiO9laQcdBSuUWks1i2qgh7lRgXnHYk8ekiE8R
eDkxj7kDxJe0mqXcceQeQtAWNPDt/7vw9hEQ02ltmfwgcbbwH/S0NJo/E+LRmll5yf0zEGSaBaQ0
vOw6QvMw8uvhT5vc3ZQOcL0YWg5Cj/0sC5f+19ksRcxrqCBIQI7977UY1pa+bsHiQwmXpYC1aP2i
GXuoncIE1jAxXAlWZjalc9O5azQzK2pumbiwAWaZ8T66S6KKk1ssUAMjXR//VNjUwRLb8MSIpzJE
gSwBDze56+CEskU3LIG7CVW5Tu8j2B+fL81OC7//YI+r3h3fbINm8OtNDt4cWPEKeO7WsY/PORUn
+ymllyyP2IZ6sVp8OczleDYH0zQwo9JZFrnPYl5c2R/GibI/id7iHF465J0/EU1icXL2VyOFjsh0
0bEkAQCcfRRxZ6uVNBPLcmU+f6Crvz1p//REGEx8QcOTKCFeNtRf6+DZfRF2vwGHmpAXEuiFy5WM
1/m7BR9TBZlfmp9g7kzV75YNGDPg/+ogkl6Zz0dAQII+C7xoLOqzon/wtvw4H8DgpNE5ckhyvNN5
rN+i85H5nhjeEX9wRJzo4fxjIXHgCEjOtCG9IWfPQokq13wbR352d4KXS7L5OovUVu8HvZG3Ynw6
KjyYDQDA3Y4UCunVBO8TfnXCXKMxZT8SYkP+DRCRkAKM/eqCFhZk4H29obK3/ftGN9al42f7V8M4
RFNfnXyZ9xAGzmJXtkpsK1IA21aoG4Qj7S4/qhcdSO9YyepkYDr89J4WzLNJ2612fyxMAvbuYHQr
RoHk3Dls3ESbXac7ZFUpEA9JYVH+nahFNlLDXoAgEAXHUjbcbfRsg3wBs1TGcNaXCNFDR2PJ0yY6
vzLgf7HgEzZwYQb9Xoz5aKzGVgIO7tU7N+riwdE5wibk+46I1/HtnFU5BdTBR5D6Y7Np+ut2dAnJ
AspK6quggr7nceQvDBeQAZa+Zy0l6dRAGYQiBVLdH9NuZ9NQNcXK2dflB7ius6XtNpQNQIsjXdwX
kNImY5w4krF/blVRAzoNGIFWIq+10Lx4uooIKfUn5U/S4tXlXJgpvgO/bId6zlPs+2g9IreY195d
NnXM7orGVwU/TA8jneNBspP8eFu15jQiHbiGeSQjdqnmrHvL6VMxNM5Y0Wgnmpuc6ZKEwuUQWyhy
M94fchNEn0u9R6qoTIUqwE6ABQbk8v0nIi5SrqYg40CdamwZqcV1SM2fic4AlRWPrvgHM23rZ6nl
G0uhfwNX9a+eN2t4+mNvOHqzzF4suiC05r7Mi3jGHTCkxph5k//hieRKT9GkACAZwPjztF3UrbRR
9R7BPYpPVeuI+Bizd2/dWHPGdNdYKpexgksSgGegyIrjFsbNzZVs6F5M3vpfkj+QcHQzmQ1bJn2h
gyZO6CY8R1m41j3aapwiJw4eLSkBGMOP9Ixq60JlgbSya5A9qnncvbg13Jh7LJ7bCCJXP4hvfZdE
VjqxuOc3A+wxF0Mfm6H+2HJW4eDVa8U/AdlnLBrOQCguNZb3khObbr49A/3XzX1BIQV0XCgA6srX
fjgC55ZV56woXkf3npWBKYpysMlVLj85wBvvfIDB1/O8g7l9xLN5Pea/2WhMvjF0wuYy2AobALsF
8EAjbo7dSlyzeBxh0lEOsFIAHuex0zupBRpyKekacp1d+gX1tYQLTBGIdq87ooMWe9tpSDgWPL10
qSfakQJFJ1vjf+oF1JBSZ6LTwWBsnArjAIhRpzMLUdOV3ElkbHTDmC1Pf4Py3tJUJJ9XcTysaZat
BWC4Fswuef6seq9sGXKX8nvPtMtRZz4YJzLuZBGo/MtHxK7p8jkRA/+0M9bucqBenm279c8Vh8cW
kQZPebWz5wXOV5rxkm/bf09Pnk63FZ1/+n8/cJSmTmic4JKY2YmDdQU6uH9kQnSOiq6l3v1X8CEJ
0TlsSm5H4HLruWyuNwuzD6kuOXqC9BNSh5t7HRXymx1vl/cy0QwWEmqsRGIbpUvAkQWfGifhPo+/
qGVRL1EYkC/Iqr8syOa7kJGablQxkbxsnG79MJ0Onyd1cAASO60R/gCztYFdhWVZwqD8tkvAyjj6
OW8HXFvAMZxN2eM9936Q66Nsb/Muyhf+Jf0FCVSADttCAoLZRmteXEv/kMGVvKqv9X1rD/MMwiOu
URXNLRmdoa/9koUk8mEfvf9lqlxsjAa8eNklLdE/bt4XIWj1JzL/Ja784jk6u49t6f4Xf0Fy2Uq9
YFVtPtiHWtURY+F9Hni9xiZ8Aa5s+ePyoOOYklXsklo6fGvRixUL/mByGUrfM1u2hjyV5OaaQx9E
OvZ+VKnaW3AqCe3Bo5V+J3kCxA5SbtxDkS5+Uxj6U65Q23Nq/mAB8LBUBjnKGrA4VuYUFnkuMLok
6Cp1zOETH/Bfygu7lso0COL8COEpi3sHb5MUM2EzQaDu0lOa9Qi+aKEc/vM1dCY0OAS+awbO+Ti0
/vs8IcDUKONEiJuPkopqXW4tELqV27zCzfLf+ytekPrftUxwnmFnMJArtjZFj6lKnLfms+Nhgyls
JpXt2IwxWVt4xk5sBK22Q4G+NFzLvUSxAISecETfN6gCCMUqao2yK+JHHjRjTrxgPBUjVebFGVB8
TFj4961ZY9eLdNeEUuei6OA6r9Hp0UfRFmMUa/7OM8KuXKoYj9jOhngv3o49A/WM3ZRTtdDPKaOh
hWt/3Tvz6yUtBCDqPoDVAFTS6/MrXn7w2WAQJyRkBP2iIibRQj5sWnh2R7bgjMrWXxTz4ull2Go2
CcqqrRGzsDkfw6hs1VVSWnmknPaJ1S/fjsKM4xykgxFDm+l1i55pgDqhuIeHmFqyrfZH8kDwlZkE
iH53wbKRM2dVIBiuqdC4zffH/EDVGI/Tap3rwdsGjXNzwS9GX8rlzf1vsR1x1oGeKivSxDUX96Cc
XhmIUHATF32K0cYzwS9tGlT5Z1GNMfmTRv7Uw+V+uzJy0AEpGy3c33S5bKx+Io84cFbGiW8RudKT
YcHUklQqjHy60uyvAjyvRo5yXFyQka3I9a6nKnTOGmsdOur08j2mtZsDkv3HrKQQjP2C380+3u0p
YGhRQxt8wDhO6FwnKsjHR3X7OTOTWKXArwORadXqF0hrXCO31ihkiA654wusm+qDBsybMiMbpanj
P5+M/UAvVejACw//rDI5IvpiS7799YWMoBxQ5dOwcfsomwysaSA5/tHTdO4iM7JpBXYJUs6HV4uD
J9Q5eIIm7z+VtKM699G+1MrOP4dK12gpNRmzHVW8iDdCDVffeAWluhPNDHHSbfY0BN8RCPSa6937
HQlNycBJdhPTAeocOuv27makhJTSinFiZ3urx6MyEAzSGuzDdn1RE4hwdPw9DsFaOQOJyoGpBwrn
pDvCxZmW6AK6xeDThjYDvCFvYkhDBehXd16gOHBeTOz4e93UzrdxUzdWiSLFtAOAiNUt57vyaVwf
nBJKYvGeoEw6zw2lUcaFhLzDfoPwfeHORTTcFYyBJ/hB+yk1RA2uGss7OlDgcurnN/4LaOOW0Mir
tthcxKb24FoWErWr6JtImtXq3RQoW4HYb8RG3N6x6eJqSAGxNOHT8F9kfc5rFo42sVyiNfQTEzcc
ysFf7CcjgAgXSMtidUVjY8Hdj3zdObJ3RZ9eoHvguebRZSCuTttBs90UboGZWdidqm6V7qN6zZhM
d8wIvW94yfMBdDxAhIgYtcJpKLXeBlFTsPAZUFsTbLOqQPTY+7zEoCE1mWQJGDAXooQq32rixHa/
MZjrRdaZTjxx9WSCxz0LOJL76T2oP6Zz8+96Ozd92P5ukMnvy0+rrxmtOnllxhp9uJGiupdxS6zR
Lr92WgmVPqA6Nvq8EVXEfMA8yM4I1sOJRV370RxC/raPEFaY1mLxygxlTGNosmp9bmww1Y09h1ST
3OuBTiWP+IAkifvdJi2xVCqRrcE5qWc61MdHCCzS7sCvTqSNcwzeRjT9UEx9tnhPbo1znNTnsIvN
Oj2/zH7iGjaMNOPFx0P4Pg9MGTcmaXh4qUzkVFYBPeZtL5gzLNkD3/F4IqMd+U6M5+rK7rEehVTP
yX9Sjpx9uKrBfKpP1Py+BRchP6FXElww7xszVWOE4yPA2ezxAlYY9aaFSqtZ0QSjLmIDeXaXfV2t
lQmbDNjZQgPztyN/ETHrWekUvH3Bw82deyGfCfEXRDDrKGq2ff9+9FpGTmDYmqIopEI4Lrnzrth/
+gRvrHUzR7/q643hGE+Cua7XV9PuYDPcqSqNSbdbeaP8fsY1DRTn++HDcVdyoZN9IXXfolD2cfW9
B7EtjZwdPDiGaXWnY53ymgVI9faCuLFIyoEOidWUsrDjQ6842NHH4Oz7h7WacceScd2aeL4uIDTh
ppoMzLsVOm8exKhSE2LnI4PJkTQHZz32tJBalDESzorB3y0+DNBWhTexp5iKh/3wJi97nmt+J2+z
iA124cgr2v0f+BIhdL7HEInc1FY8uQxCBk4DQr9TzA+eDz6peb7DpVGFOge/jh1sd8gvnlSkp6uu
AcPlZ6aSNF13CqbLLFUs9J/5z7N3yqd7qCoFIwF9yE7XyxksO1An9See+OBl2PgEvDa3AfCLDw/7
0WpanHDpS+/zpXZIVX4PJLBuNjOASvb8IFTPuPlPaYcp8ryYAzTo6uFUsR60Tsr0DlryoIGzU0iN
j6oNE4h1JUfCm6arVUC7VTRq2dW2IENX/gYd2HLCyi95tqXIp7v7CQoykZsYivOPD0pqR33/Fozg
OVfMm9V2ugFsRI4k3EP8ddz1s24BVyxYudEyrncip7LeNKAmGKVu+XW8kUwGb1fr2cul0tY7l6tL
tSku8qh+Saj1GWOulwoMbAOZCg6/NucsILJAMcqbMKkQvZyVLlGNHouj6I/JVdUR+uwJP5fuWRrj
gMn2FCKL1OJ0HHYeTFWgGAKFfjkJFaD613/4FunSDtYt987Pll8WC1tkcMplNk9XODDLVnS7JW9x
qK7A0xmNai7dBc3xsODhzKEO67t+IyYRtDWQt/Gu4gjAzffIiF3Swc7ORTATGdG21zjdepZ3b9QJ
ltPvLqz4PQMxOd//Z94ym1TB4hPGtahq3hY88tdQiZGIL75n1NqS8s3rfG6cnNozFUNdGS/C54nl
0vLWRSi2MzXi2Sl+gF3vRssc+wOA3ZRzQCTl5dn2sxo5S92RjnRm7/jjoQkM939MpF9M45sZd7xG
7M/Q2WZL51xNlifthtzbDl5QQkATBmFcN4GcP4M4MzF0k/l9EwkJHpHf4sG2Wx1Pk5YWn68nNrPZ
x8qKykd9qnYuED/pC4XuovhAY/tjKWQ1FuUF3okNtWQM3SaBTgeJXZbKE9GT8P0oYYwcPOABh1sf
w0uIJ4EjGqT4Y81dWdtvTffiaIZcPPMPcY0g3qbYh9ABvvytAG3ZGXTFGB034dopQ4irtWGY3xE1
V70KcZX6uUCovmZNwYUzB+x9Ce0Dd2LDr/5k7MUGGBkNqmdOZEc5pXc0F8tgZDyR3/vBrxn4hyjW
NL4Rvg+hhYbVNaTn3LPvl+svOoCu1ONWLK9248Wm6HVSGxclOte8lCF8HSHJp7aSu3XEshIDVEx1
L2EtxMAuw043p4gA8M76VExDJu0My+QX6diXxs7a+sYarm2kcFAzhMvMttRwORtUPmhobCpARWnS
iaBtMSELH2RMA5reo7Te/TwWA/lJuQMC9qCfPKJj2v+4+g1P7o2VB/3grT/9Dtpypmw3hKXvXTda
mBMVpqbsf5iWLPzkHNYFRIeNyC3c4uV2/Oder9s1X4O9Y3ckyoRRaBWk1DMUSMO4ajKaiWATHjOh
vzRt1PqKAvJwGH0ItyT5X7OJhh7YbRNTwPaDWPSDEFkOUfc5kTAGYibjJKHSK6WDhhzIzaLXBl+g
dJSuj7Eqt90HiuiRFWmL+OaJ2l6eUO2QjTjgvhNF7Qszdn0jKhTyxcbkZDShe3FYR8+w50SZg6y6
+JrKSCYQEXvlmxoRuXVHg9oW2NO7N07p6hjWNFKBnunaNVOQ1NddwMiWlMpdoTrf9A/Z77W7Sjow
9uo/SmHVcLphk7lqSm1yHKyKr48zAVEwggvl2740KRkOTHMQU9wgDvSNKz+YGhsZkGeYOGvwI69x
5CuD8zD1mcdljrC4r3I8cJoEZeFNYu7F+RAbn6RLZBqLXGGSIoHOrLaGmZlGXMrY/JfKbhFtjYaP
i6tI+mVsr1IL7hrUYXk2JCIPUiPEQ3EmDk76y1kIiKYOk0MQvUkq3hgXt+WsJbMG6l7DOq0BRNMK
iLclWfjHn8IbA6nCAKLhq7r90zKb/dhxVg79P2+VGjoybvghgBbyOEMRkik1D52KXCEbamx0gIwJ
TrHD/7i1n2M4Y99Vk9eZL6eyyEDHYRNfZixsg7y/JSOWoaiaytX2NF+/UDqUKI8OIN3xlXA5GKFL
EFHi6NMWeEmoy4Sw7yWXkZkd0QaEpx9N4wuqC5N/jE2vIONM079tjORhORPkpYEvcFAsWbO+sut1
kChGRCdXw+nmGcQ+vxVHOm62+IcX4j2uhKctvShu8/AGG84IOhPFj4bb+64T6xJ2WXDxtBmk4Ob3
OTIwu8LBOncG+Fo5mLsqyX824cQHPbrWwOleR5zwgVKhL2J3wk9t226Zjs1Af8jGOYajhm08mfwJ
IvPAJAuo4+EB/fSBwkQ4LRp2JYdOZbWu+lXZtk+iMpXRWB3xaflDoacvGR18+75SGTOfp/1RBEnr
phFP/9kMeE889C8BrNIRAbHmjv50Ub1X5IE7XlfkKUE+oEFjqXdTS/LJy6YdpJgpHC9goadondEA
vNQR17kyKmuskXNLnsYJTssj23Tt0srDinfJbnwuCNxiGhiGVlfr42MC1Yn1IDVIRd3Mchggpt6O
+0p+8fa1e1qhUwqOBdgZcoVP8p06IM3o4d/GDX8HercLM5nBMByTBZEiHlFcqEE9tAUspcozClsF
aUdJHVsoqnTbDngNjk9kkVn/k42ks9ofP8H2DIsNYtJ1i/9XZhpDR44enCjh312f82JOhhmh/alk
W62nsL7ukCss2i5TY+Oxt651XJWPIp349lZy7aq1Nd1sDIoJEBkAArDM3mZPlTOnCo08QderT0Nb
4jgPbee8uSj1qY34DQB+nmiBve+QiRALpAiXUbKBwXOmsFQmkV98OQG68s0FErKAVPStSvLK1C8k
kAK5zxxW9tkvlstWaBw1/Srf35AcpSCB5JcIx14gbxlI6jjA5Brgt1xWpuwdeLiNiL5+EuHVfO5M
hP7Ruj4oM/tMYWtjtCk/rVod2sQdsHH73N7un8ej/zf27GMtoOgQ4BTWdc7/iSizei7Qb7KKQoa6
HqeavZINFR5ytS/1VCTmc5E2jIj9g4nGP73Sc3Sd7WqYR3id5mzcywgnRsa5dXsgLObYDpfbStlZ
89gma9LltbN98rutPipSG+VVCZ7wESJRs5kIPSbz2QvPeyExS+FCVXtL8/C8V+jIpfmvAr25tFCi
P6bbupJFUX7A15hfIrIOMi3ZBKKdQVwIbtWH1zb1W2Y6HPznf75gECv74sztORtCWd6tyBPwnL+O
xJRFHSg83Y2wxUehixyWlto7TZ45Zl3EHohZF1kSeY1iOFPFSvYLF6+2iRIpZHDvlz8d0VPwC3cK
ewb65Um5SE1KTJNaIsHSqmm9YRssTo9FeHebdpjOB23Iv4rgEC2JiB48Btgj9VoRvH+zDrfyHWJQ
9gmrB4B0/3NRO9LTORRRAAsvhdOytqvGmn7FOGEjQn3pZzTNZAzfkMFPrfOnBESmT+WpnBTqWIXg
7ThTSMDYN60df01XSxwQydlMKVGYr0gMoEA/HTXZqTaPjv9ixJPP393KcQSs+WFLTBys2VgIvZE2
JMV1OzuFXpSxc0oEVGBkPEwAZWpYxSQFFqT1I4ml6ccQftQIXF3/eFfMEnV1I8qGswTlc9WrnYR7
/4Hi6DOzQ6NXagJS/EkpXax5fuPfhm+7hqFjMJlA7xuiDWRr9mlZLpuCZF/QHfyE0atuQgAjcscO
D3M05sLsWlWkApie0IYEJmvEBXjgzG6W4opj03yn7VBNItbSxy5g9x6DtKa/TzU+T8+yFLAYfpsF
TLeKpCjE2YxMavGaQdRA1yiil3LW0nYLRTMgsh1YvQdAvScFXgbeFTksl4C4KFE7J1SYlVA4vOzU
poIXZWdRDGSSW+tD0av47GLZ+ms5Lp9OPIoSquC5rrdx9UAS2egWo909nXGxErJx5HLTru/WzNp1
svsPZctcfBckUVbJd10SmVTGL9b02j0S5gvkRz+v+fPJA5Q8OR7hJmlTZsrToRlns650rh2Esoag
Fy2xUcj8QxFkZooGNeuurY+npaWbW9zQ8ZnfL65Q74dFaif3NOwu0gq8ipoXRJwvqJyxq0HKjYy0
s5RRhIf01LMhabbPOlAEhJUID1SgaOxEcjr25dBqeki/mH8N835msxkmT45eG8RwjohD8XbhS+Jt
pQV8wVHwMIDonlAtKXxz7fYmJtvz5/sFs7oTU7E+GyTW1joJUS6zNoKYnAt0+ijCerYMjZooGaDQ
KxXUmszbU1aZWodSuCFfMsP7lROVWROYSqoKc/suQRbrsehbkBnYH0Rg/693SJOR3YwQn73hcxpy
PeXyhdey1m9pMumUhhtiXV3cU7XQG0dQF8ldA2TrJ+ud9m8qyRsXMQLQMkW7QAQ2YAfTu321BNXz
IFhiui0+N2lrFwrYFO+KxRfDybhg9owR4CbXM6DiBSSRvJ5ngDnyn0a36GZpiblZEZhTMWGJGANB
TPoJwnwvnGW3+HuRWNUsgxqvj2vcRSVUWNEO1iNYkRUON9IMq/H/yseZbHHFyWaO43Guwm2CzhPv
Gq21s9pZYuUJtMgc/eM13Ox/tvUS7zscSly8E2CYfp/DTIDz+OlRfeoKW7PhH4/Z22fshi9iHM+N
WhBVv43dpdXe/+NO2rbj4qNzri3nESa3fX2OcAd6wXFr2zP5LfuU823sMmkgjD9h/bogzJyvX1Mw
PXzFeXFK/vMN7oaha5cLw+hsZ9HqVjlp8FpBM0ZDNffzRPszt8trUkBhY2B/cM0YPHE6mce4bjks
+5zo210HDtzG54ehI5IRxYyFiIWMVnaS1QWL9XuljQlpVwbfL65Z/jzgpwH4kKdtt2S+KOK1HftN
VIBI+L5xGoNmkXgdwZqXLtAP8A0eDVGM6MGmbVp9+uzLVuOyeEJMhpHDBDQF9XCh3gVQMq0/kyCg
qmK+DaJddJ7YRSMkppSw+fFCIySvvNqKYw9jWyOiAs6O6/MCqIdzEfeCuABWDyjZzrmZOy4sKwMb
+jOWqcZPjj8kEYYJMI1D3/gtfzb6wRo/b4wNk59ShS+MRLmJJuBYIO1aT0n5nfr7Xs4n1eDqSqQf
/AWbNMCJBxFlJ6D+f/OR8cxNgMC5ld0P85Jv+hstwo+6EYM2wRNwvib+3/+NOapFcnzUIVaGUWHw
BHN7X5X/LSgE6ivtNwtnDH2Qrbz9NLp/eG3s80OzCZ1yeCZefgucgwxqtFrbR4/igN5I5FRWWeD7
/fNdxzM5ZHE9Gf3f9VxnpjB/9OYohApbx2HIAi7EraNvTsLYx6elV0IsArQgDDujKRg/OaFNg4lv
PgqSALIzLAw5ZVGsKPAUWDXlFL8mPWnpte6E5/OcRVD2PYnHb5kGzQAva28zc6fbmUH/bQqH+6a2
BKFvefwl/yXiskE6vNXCLloVbqncJdGZQa1QtPnOsGm2Q0gB/Of5uVr891oprfg42PHhnOusmDdY
M9Hq4st9DApkeeT7xn+Q7chIgAsZko3swvWJb5E48w8kkARXqg9t1tSv94dEJeaQU+CJDm+h4ndE
9BDDuBjp8dUTHH7RnfU6tMZqUz6P7AVcRiXBM5GIrayQ/QyQg9tc2KvfhTO0imcMT/YH38F+CDvh
sPUJw6vYr+Ytyb4AJ9zHCt6vtqXp6BHHwKlJEdeyG9pUSURo7/tHED5Ru9b66cf4yoSHZXHiB2pg
RQnq3TiJ37jliMaj0obX9tVpFYILl4c1NJEAI995LLKct3FPMIqemNDVa1pp9f0JW63SjKOeP0Zi
yj5jjkgwaY7wTp0MZniWJm8vL2ggGt2mkBLodYfOrePYy4h+VPDZ8gEyoQoJVRZwoK8dsvVlkKAC
0lrOGHjOd5TjCyp2FwQrN2xaDmmSdbdM8L9UEu+9mhLkZuRZfiuiffZJOzsHjE3dXiu3HjxM6bCe
uVSZ40Sh8yI6dl/yQaeWs2xzSNvYZS6nYx5IUvndVTBhDVHfQ066QTF42qeOEjbWIFWF62xj5kJp
MhWBpQ6oF4Y/4IgR/16yHh+1UEVwuTl181gdwvjCIdiM7jWkQ/38AOueU+KKyVW1NXM8Oz1UxMfe
IvD6vRfLhObiGYqq67HNkQEhGA3hN35bb3d8Y0lEwhastITaTjWtjg3tpUyaV3SGvwshKBCoOaYk
xFhJEF2RfszzNwkcYOTGRgqainPzslF0BesitGMxMmefv1xKxnyEPATbMvr8ynJ/cKXWHavIxIMm
4ceqYLrwaH9g5t2D5W4RKCjysCxlAEB8Jo0o4OvdsCM3+egv2y7wqA5SP6q91HZhXc9X2eMWX9LE
/xC4VbcBe9O02WimoH7NKzDXx9wOPxkAB3jYwtL1sTuZbuW4iQ9qFjXP/hm0ZJLRm0tttOt2auRk
IAckfbWXAellrGl4pBNrffxlnFQp6sA177S4rZYa0Xsqs0KMYwUa2wxO5tpSQ1YhXdgP86cvOoX9
RFSjOPLUlJ0WqnzO9qzpOPYxlPc0UOva0XTl+Hx2wPXbmzEsEfaIdujeGY6qaZI+2lUWQ8ik1OF6
CBO2RrB6vWsdVVbsDTf+uQDdEQQw9vova0hGDm5gBG2i8QViv/FCFVYpXhdejtlEWdZdUURY1QvP
1LtQqKSz5lTF5+3Zn0CSQb4IJpKKQRRivIAe9ie5P1eSy5qySycmFofl2AlMmlQeuR/abm4VNbj4
RgsxVY3jVZSSYDBpiCOL5fI1S7eFFUcdrumSjm9O55MwoALdAnlvdZcG1sYDLgfDkuzRkPuJdzOO
exT/JAtp4msKFj1KoYA3RJp7U5CSffNCBYwNAa+liibVTNIJXOuRoBYsSjhCmcb5hZvZBOucI6Nm
z2n4Ps0Ns9N93Vy4jjBBXV7OZV3pQ29HR6I2GO1+3H26ANpXlZhtaThcLCuYFFkqna5hfoDE2zXr
b3NHcOOa8g+gBsukdfsft9kLlN1O9P0GGk3fAeHJOYBAd0ZUTCecl1kTWQCN6yT9YALBN+bru7VI
fkrfKFYfxfiRrZBkRjnAQiYKAOobeokrfEFAIKjcxE8X/FFMBv8gs20s93FjZja0ERibAQ0LZkhW
cdv6v8k6LAUkZz9gwHFPPbsYvOevjyselYqciisnUP2c3GkmnQ41Q2Sscqcp7zU+UvBQMo43s3JQ
mRMNgOoN25iPdQ/x6taJ6Z1STEwfT+peBJX6V9uRvvh/jeXf4k56ZeIyb7mFFYP9zFaoEdkvmVQQ
lGZDpUWiXLoXyliIeLhKrxjDtDqu7j8zUwI/b2NhYKjUdRYOd9MwcfFyIBHYwq7sWtpt07a++BZe
FNEZRQ8wGNxoPcHBT9v8qEesyp7w34kjRA5ySkNFpTEcPXGowh77x/eRChO7qhwxs2ATrM4Y8wEQ
crQ2wxMmA4kC6NyYQMkYio/iL25vvuo//lwA5NMh/+p3Ctfqfr4dUA3aO8+hbWXjAA8uupsdDvIH
EVgL/vm5j6txADWOR3jBWNastTSy42XFWgXWrMHbGZI1UcixDoyeFeFSyIihCDASAveDkJRnXoIQ
lhDNtcU3u+IFFED7nbXInaAnprcz3vc7p3IghDQ0q01GrhrLAqc1Wora/HgwY7Khd6AgSi+5+WXp
AQw11WXLmHr7i7Hcga3C8vn4soREnumn1unyYiRK7yGGQqqAQX0CahfwhHiXOjSGgkk6j1b1iEhD
RyPzLcD2ru8vCEjQo1NYRBOqotjgLIolFSi1GJnKFZ/V2rX72tU+wJ6T6GIccHDE/tP9FaaQVv9i
k7oucdW4LytUsccvFI+6wjY+v+ozurVX0hKG7IuptZARSYQr0ToVkueGhP2MAycGBKdTAFFMV+Js
0UEJ3ApZiBCicOepYa9G21nQBIGdiKfAB5LAblTrn4sf/zEEK/ZCTRrQu8x72zCkCaumHHEnb2YT
bhmDQv5x2hzFudR6ZjV34OurZITKtSBrW75wO4yJbYIcI3EG5dVjqI3gq0CYy4133yeNUSVb4fKV
DK5Y0BQSwcwGT7i0QVFMnP7RDb3HWWAJevbpdy7QJ5o26w94bXGXFZBA5s18CsDawh1LRrOnzCda
z6SRgy71hcgONHs2UB3PjxrGqyoHL4BoydCPTBev41GFaKbyIPuz/E9/pztpRlBBAYCi3/kwRHma
j3USuywP4o6eClHKXNeh8sXn8wMkeUFB5SX/TINUMDS7d98C5nv6qrGkRqSC8T23fSAeSIQOjF9l
dgF4pN8rIpS9g+1FclUsxlLqO/gTQR0xvb1Sd3ioABvTopjM2PenudAWs4vNPRruqxNBilxQTldN
I6/VFSVemyS5yj2GOCWMTU7kgnJxea31onmFHh0PmDTmesLD3BK2dLQDwQfsM61k2xB/9O1v7VcS
XyU6jUiByn17eBOpLnAtd1qFzwkXGunQwwunEqCkAHelP56P7WJXtwxpdDan9/q3WI8zT67icJlO
HvS0ikyfwWrTPbLU85BkIjfYpyltxR+xykqvL5DR0ozVYxdW2c28d/ja+HloXN2TU+uXWcE2NUY9
bkYxXgUtFRE2g47zEjjKFO5H1AVKojgWdLYuV3QmUWEGdTxNEmqb3V02w7l+0SM8282tTVmkO8ow
ZcOxSwhArWEoubigeJ88taq/7bqywptN7zXAzUBFV5XnqjvGy6WhkcVcGEm5TFAJ/NJ9bHMSeRwR
MK2/ObzFL0w5rbLU9QRUwN5ZdEnHRyL58i7x3RYLF7JACGY8JX6qDKIcud1VC8MaQ6bpEtJKeKeX
ZcIAO1JqDgfblfdbhJoUJCNYx1RSqxsxmwRMgMrYJgK+dEXVrhPO8/gifeE2sz7aU7EGe96Axbyf
rJptRfGgXlwQoBOSVtWssse7CuboBH0sPzQllSCp3P9c0QtBTQsJQ64cLd1X/jZFEZf5V2QPz8Br
91L2VqX7HCSD4A6LG6T7nc+A5MAvjjry2/OytezmVEAlxMnVCW1Hmt2tDShIYzOLLwaC+A7NXYJ2
k9uOWy+6NVknFYdY+JfFXKV88uKhLGWdWAZpt5gFYJHggpbR55fBp4juJGd07JR4dIRo1CsZ5dUn
sZ0K1vNdtSUISeMYQJzvgkajK1+Y3oSShgsd+ClLNsPKNyQq2djsr2bJRpnbPazu3Yfo5yeQ5nEf
00QgsFZnE6Nj1X9ZTCKyW3bajHsWFUs+Sbz1K9DwgfmpO1o5qvTeupJPCVbcOCnAZL6dIgIWwSdm
+cwZmtoodcaUr5ry1CqsfQL/cW1oZhzruHtpsXG32xmfNhdKuOhLOct3OCp8xb7F6qjiqNEZh7kp
dD8lSRkFFuREbxQmP7rzx+uhzmdnofy5Y06qOnCPzYfqrPEIKzu4dNXZxMxqJQ4texg1F5KXSkU3
zZ8iTjW79CxfOaBVKGftLJdFm8HGz3TygVSz7wnpWPihIk3f7vahuIfmbzSjTjmByV28g+ym5JfD
QeZqRaOHcbM+EAD+RebfcGjTnPierajwOZezGkR0QAM4Gx1nDnvcNhj+PQutq05IGMEYjZSEOrVX
ncYii34zAu0DfrxC9eB0fYhoJ0xCPnG3JcQtaZBRzwDhbDKowh66jY4wvRXL9XKe4RI0mb5S5/Qc
YOzdrQw+ebA7rymCaKhzyjB1FjA2ez12Kt1OOJ9cLOC+JhDEhlaOTPk5OtBBhEKPniAO5ZZV8Nwz
/O7vzi0BSQob6/yPOlZW6sP43CLvSW+P7QlWHOH/SiXP2nfJDX9dZD1jO4MxH+fLWfhoTwVOYCZH
l4FNf9jbRKpsiqmYFXL6tXkJu5BF9ybviBT2TzFUPBTbHyBIkGCtnxN6NYJ4d5a/RUpkHhd4AEvg
71Ou4bcabY7HhozUKaDWTI3R+5DESUplUHS4E5TnblRaU6fnUusN4sM6NSqRbZLw7ggvmMzqJ9y7
Z/OegHBHKFRdV8GdBPkAdmtNPmjNzAx3nLNnzVCR0jW3DwwJArkoR2N5ki8onmVvRQMyh4fVkePJ
c1t7DVNWYmHUwfd0DJBacmxcWOGN7o3uNmFQNpAVNhd1eA0BsT0ODRndnCf9+iuyi1Ja2gzuO/N6
oPrnWlqia3APLkY74mduBOkP9XeQPCpw3mwBZoP9MEg6g50xJW8z/8Ei5efV6XFR5xLpyc/cyjjM
lvKiEkY3UrTczBXpK9HimCR0ght8i9ZK1zw8LVXmkk0FHCxbQ1DPybyqrBhg165W58rVlZ/CP0Bp
wIIKYI/zvX7KZcaXmouJJPlrvcRFAcHpEEyUfBs43pObZuQ6f9wV9aMAy6EhxhmGsNB/fUU2mkN5
0YsQsY2iyUclvOJjvoX2wiQdzsSorRtJK5GUrxzxgcjrjnPte1mod0OTCabaWVi4LTNTev/vk/I2
XmyA3GNOyzgOt1D8i3BMMcNtH3e8AXqp1Qky5oXv7G22cdCr+iZJHnX+2qpdTHlD80xSe8WO/JUG
QgR2WbmQNLvU8nkPsvNVW+u7EF0sXgo+LRMbLtTx5NB32RIr4vauBP0MIiXATUlRc86bFqwx6Rit
8j36Ob+C6mQgvptqXcC2VhFD2AzHW2FqIz6RYsIYAKz5YsGIHjT2u938Vkw36bB9r0bRB5nd6qgl
Ing+l9Y0Z54kYYI7MvtAbSM5RUJfrPzqwXy0DbzyWHof5p7ysmF2j592+QP5998ZqqKADnNKF1Wy
rIzclbpjefzyELgTSTTsvPNDDOsLGX/xivb0Qivos0T/DAE0fNmjCxvKoplOMmanbswC13lucJw8
U/8ED4tSzoo630A6Sh85taQJ4QMCAsSNp3W+Bi2QuW8i4BFg2huTYPhZQzkDNRSQ669lN8bEqlYZ
okBh3pU09UKEMh+hq/GHBWJ0DG6lijawxB1Kr3/t8Fbe//Q/f11lHsqfuJEW6KL1A/TkErS48669
vLmZ1x4HM9+/GnQEC4+vpDuDQLGJ08jVw+gUswjkGcjQfW6xAJfZfYC4Mw/ujxa2IGNb4owgzTMS
yBb6qMokxUHlMJ55nEXJ6H6816HWsPLlBgK8DkwUPbPrlGvbksunpkZ4rrSwSpEmTibsdh0+pLDs
bsnhzrFSMrY/41tQXNZYFzuJirnv7h7OZ9o4JWFQuhvXcH/hzorMOjNsVp6SWSGHjikBv0RyswXB
KWv+8Kquh9SMcBUEIDmVzd2kS9TMmyg6ISdHec0UrUngtWBGdvCKO3EiAclp+ztauRo9qBK+00nB
eaihLyVyFBYxpQ/4pIXcgOysVWNV+ovQHCRIuhbcHQui081+WR4Yh8hMyjM6qtED5untUDf/hLBJ
1Ur66P6xbNgqxWBcL4seu919it0fzcd8plDiemvx8z/pBGwt8/ssmLUQi0wjxS6Joou1pSHT8KW6
tG5QVt0iofmKugppHuaivgn62zZwpO5teivEhYx8xrCkzLzmdGMegb72K3F1GboMpu7HZ8JKFUJJ
3yqdhuQuDWuSEOOkRDZqXHixBKvGKDZTi9MYXoWTnL5Qgn507MYlQQelwvIR0mBSUWFRgTQb8z+H
oGD7jvT1fn6Uf2loO+GZN46BOylMTB9LKmwYvP3cyEHurOzJusCT446omVWrxOAeLEiDYMrcE2Bm
nNYakOL765pK9zROZjYlb9ij2gTwEEH11Ri/l13ouwxLlE4QawuJAZzQTwIbyrQNC01ynXfGNAlu
IBPBy7nwCfR4OuXJKE6DCzpr2QcmoS+/uSGZauXNheFjWVnR+1QnFkKHN+tqX6EGAneZm2mUxvyl
XjP2nMyW0qAmupyCwpHbv1gHuMhC2PVqOM73Ijd8Dk2gzTyB8r9I5rYr7k8WCyTbJFxjLnIAnH49
0AxCRieEKQGmgJITQljpVZJqvuTYqbuBeBW7nl9QAfknp8BZwnsfTKPDrm0e4iNZbfo5xkUd9Jtz
8wxdIUhnqM2qsP6tIRrREkY24voi51Ck45OqbF5HtJw/IqsK7nCiFOcws/x7Hxmsu/NbZBVlSg2z
pp3DbKqUU23QfvGqMIonemqAlkBSNEs89u1Rzj8LfNK79pg2PHwl0DYE0FG4YdP+0tbtvR6PNxcL
lIgtfOnhWD/eBbflZfwoO5U3QChNGWYfqR01ONc8BD2KQ2UykWQu5NwNlk/7kOgvv34oCDCwdnav
KKgtmmHh1gwuxIwvFbHrmknElW5JZ3pfcolcPDKhWxLweLJAKE0a3Xhf3a73Bf45A7BGpsYmt3eC
YgViq4E4YNl0oZFZm1lWqw9dJCuUGuatNBnEn8PSMjHUDa7w17Kt/u0brU5oOUXc/6jLeqm7HB91
djUJCIk2Xb3GzOEb9plLUQdPfvveUtLdBQZQk6UqkeMAGD6d+aLliaZBXVLWwC0Yq15/pNVYZQrB
GOE+P4F1jJF+34Nwm2H6WPSOFecBuz2Zo+JQxosuom/eIi7uuH518TetOSdW+ZXtzUVZHBrZkiiW
r/dAKvw5H1Yksnq/4PG4gtvVunoL0hJ1CHn2w5epD4CSuanClhEZMvK9OMP8AAICja9yFhed92zB
ROhqeKijw8t97fsupCRtd63K/W7Ig2AaXiDsqqLs3JggZPn4LiHzkgTtd25sOLQxmS4h8sctq5yZ
nQfLctEDtx8fW1uR9inoHRFcupj8BE/a90hDIPPUtOQ9nhWyu3ig8kaOMPzPk2Qy/ufZsxdfeqs/
ehXmEZJ7toLXSupXZw357hwN7lS4RU1RgODpymO4JWhZuamnWV+2O77dEqUyvNOGjiXZ1JA6dqO6
H908tvDem80gL66j+DDiY8SpCXhK6OL7l6MmVcPxLDcSC8Q0/GQs6YBrkFCYxo1fGK472mRiXTWb
scEw/kOOrDD8nyPq1ThrWruJScA2q40SqrCZLA3Z+WSm+T3nztNX03va3cuYZOSywwc7NiOa10Jv
RWzcDE4L+YdXqipYRiIiKNx1fxH85etpLYQ5fu5Tv4Kv7N4bTs78NDXlHvnBBDNr6LLp8KYt0PFJ
WFnH8tvL0PpsSB4rPaYS+oK9+4qGxkCsZ8QiM7rsNRSfoeL8jDrJ/Kv+ETzeSUw20VQXMMR3OLro
uKBv9EwaiIn4KdLqe53MY03KamWtUaxhii6Ibzn6CW55P7pkSUKOLZcd3d1ReHmzKmJ7B5Igt/YK
nJIJByS7p+FeBOibSOuJ3lLgqD4HNEYmnSfLtGmG6Etlkr6VhKW+oTtXt+kM9zcjTF26D35sSyKZ
OXOp6KUbdWoNwnydXyx+SqTKwTt2fyDAMqq/51Jws+vFGlVpelJyT1MlUI1xzUnuuSNCQyqlb08g
rEH/E0noLZ+TELgt+J/0lxGqfJpa0uXm8c0nnbLIyAxEHMnuIPwW9Xv8fC4fIyaPrn5VhI1aD+IG
WsKwuhvxZALooAZ775mN5heZ3OybExWuLbEaie53YYKtFapeOEKwlC96A1bdoMSApGfeXf8eekeW
JaJ2U+hGwjiTgvN8mekO4/5tu1dhNOcQDedmAo7pZbpkH/aSu7LfyI8n0eveoDZV7GcxRTG5QxFK
cIwrfEgVdZvI8NoZTUQ47mo8sKBCj83hCH/dMTmB1BAhm2oArMd5T4YG453siNOh/bh7ynShVX8m
7vS6Y4kPJt6d9MDpQZQfjSqyJGUshhOQwvoO8u7x5mvELGxXfwdzLnH3vaAwoCQdPCRxatiEZwqP
BWWTdQTdwDE+53nCU7wm+UxzU57whD0F9xmvbijhbuxo5EoM8DUCFXjwei7A/N/ZOuhkkikeNXvX
DEkEgAOPN/Z80xeA2Tzc+XjQLuRpgr2KhmLo1uAJWhY1NESv22IAVYFJ5HxjkrMcqpGMYGYCY34F
NE0P/COTZa6dLGBGc81ekT0bRcWiQSKGajDz+0JpP0bkhURBvbH/e71uNnoHanxThALyb1NENGeX
PB2gPBeTXgWcwTA2joD0uondyOdw64l5UR203PepQ1gSmpsrvVCj+hQY3skWvNuT/q5i7I5kN2qr
XCAiovLjbvd2C20oK+ExvddSSoC0av/4AT4tdIv2sHBSE9Q+n4UEVAzrfr1Szk3LRqxFJA/SuxFA
I+6AgDn7CSb80Lfyyr+ERwq1YMpTHqY+TmT2yomRaG0YCZd0jJinNdbFN6H6YsMlFFxZ2A8/ekbF
vePcbQ05nuK16+tDwng491TXx0GmauemA8iquKdz9Y+E+wi1f8M+XiFy/6NMaMGOuvX5wk8Eqm9C
G0eRYfLQxooYZj84TCu6idReagH/in8GkeRLPimd/Pndh1fd/ZQNO27IfPGOWwol7cP7kfW2YSdR
pRjw4v3MekaxRv7JVmE99/Qo8ENmNcm4N2UxWs43urZqReApilcWjA/gi39TKIheOpMI+qp7lz3T
Skh9Cz5w+TUB39Kc6ZpFWLbbqmPK1QzKEbWOAoHYTdMkmt/Meu6ed8Ef8N7S4cSRLsM6s3AoufJC
oDuhx8xnmY5hTvC9URC4iPoRdMVHji/y7DQ+VjN1gklIDwhcJlrTDLVAeRL6WkvEJyDBtuWgfWxi
LXNC3Zpniq4ELSjRh9H05tQQDK+ZpWM7qaZtvhsb1rDDhVSos0k1u63AhkA2rakDySGdKMuTUeFJ
8pGyFmTmYYpBqQigKT3LnvWQpLBjE7OEwa07IHqtunHfBXvugOKHItL0W5p/FIvcU3PfvCe392rt
Ak2sQCEJmefHgLU95OREP2tFPWTG36cugWcop09VKxOCZlkm/0G2+NReRjmhERjIMfYs0pBsy9NE
kfaeA3N6o2BMWoCxbUdLgZ+54UrnFhscgLD9l/yvancgyx+doDOBPsCRGODBdmM96rQYuTxxLPFK
z/AWE9/TEFoshofJxmwcRfJxABSBHitMYzqB39lxn8pXN2252CkVVqPvSFFGSHMXMYt8hdoR5Fo0
t6LHsCEiQi9YJrybVb2RCGYEuvaFImkGvFMHL8fxMUzB/3gQOXjFUSTzqb7ex4xqR4bBTj6kqO8Y
akQcmR33GVl13EsqCMMH6UoTpI+rjQe5VnqcdySyYvM1u6PFH1O9fzjCTKMxRT8YavvvB2P0obYb
JgMLQ7BhjwQvdEOan7aLa79hGBd2d6+QZqJuhbHbv/T2uzQy0gKmIzoNDDdmhHa5CvJ7oDP11JXl
WE+GE0mqx/rAuofyKOLPZ13mVIMLDDb5y/0qQvtm9m7LtsRSKJKOVCAK+RjmHRa4nyXAH5zFgocN
mSbDW/OLGgpdmbUAwuQ0JLLgstBtChuDDOV8C0xp6V/Q1tfLbc9LOC1kjKiGFtTTs9l1PfnHQgXo
O7s/nj2v7Zz69eHMyLq7wpFaUKLhkdv0hO8VX699A+NA0ZFmeMSLOtwngenuCeHt2LRfDulWjZ2M
fIY8QM9AjNBHkodE/TfbIkChUgMvN5T+xNecshgUevb4NDVml77da+N4KGhUyjqJlI7RkFN9DTF5
QCgkZs/YfA6uAurkwZmySogKpe4glb7fxbIezlayadwii/jzBCdkBZZ/4lMZoPLWwLNZrJ70MnPD
cqa7Ou6wURZbxnqxUAY96niw2pxwc1YqjPQOMfsQvXukiJasqHLakWIMuePl293T1uKNpTUSW0Ty
9RwwfAgmtZecNXgrlHsjVUm0963PXYbbfPYH1syLFXyrbDOa+TL6DVn50w0WlJLY21/L+8SJEERK
gCDeuy1OqkTCHyDjkMgZ7ibwTtmUHEid5HhTZl/wnsfVEIQj8mHlP6C/P8ncQz1M+KgqA6eVsH8h
iMnpc16Ulp15nZu4VocHD2up5ipNSl+MIMsYD1VIL+jlJKNbtq7eV6vp6D6HYd1PZ3ThKCu97XIQ
olLtFtSYVF94WmRPE/Mz+/GZUid2ti55N3a25U08EX+IfLgS0IM9JU/ZyltU/QJ0OiWwt0ExLpuR
7vRerjBGQZSkVcR/rr1Kp4Qwvx8aq2YsbM9ZvYFGLOiqPdWhCjTcuVet7O/2BMKuifAWw2+11mEG
4Jkr5+/v/vy0p0yayBpnVYgDwDybhoMYA5F3lJJXVhO5GU3OvymG0QdeoKL4FGuVwFPJqM2DdPyk
1vvraeKSqThr6nAzH95GwfChw5USjBcFh/y5qXWzsaFMHiDACh6cLXnJMqw9+5tHohGJ8CwrD7Cr
lo02SDItBSFtERBjXAOudoeeaDNJF87gCpIL+mUAm8SqxwBIk35fndgX23hnUb8NQ20MCEsqLVe5
dES3IcafwMmBfy9OR7Pyr38xoIgNYUnRRnG1JVYGVAjqkzO4lN6uK6RbjR3xyjc6D5WPGgESdMFc
LefOjEeUUWTWpSHGUgabKoHhMubGFZwxy2vhF4nuxYNjD0ZbSsd2scwbholWz4DnTqdH/UAa9wcV
uLpfObMo0o6/lXUoEk/xn4MOOk3J19hHezG0c9hhTFAyRNmJM65Cvr4dRg0gXECwTKj/w+HwzFQr
RkABttya0x9bQ9ZhzRlRBRCv5xy/c5VVg3Wulp3KscL6VcRuBXszs+n6UfaMC9YKNq2y2a6QugUg
Nt83vIfObI4r7QH4aPpQLXqqN0jz2k7Xa/xg0cwcDxqkzXvKHvTQIhq2+Xn4g6rz+DSXqTqtlVEm
7pSQdq8ZyPh5m6tePR5lSKSe7OJ8whljSeE+dPz1bUh8vXBFh0bVXgfO1iBnRFu1T4ELm86nX1V8
d3fQ0A+M5e3YjR0pGNLl4/Wy68rvawFhQ8X2tB6mz3HHoYng4XXUSM93JsF7yJGhBxQG4eBBZnMd
LUIcm8iCYqTQ7Rw8Ci0XcYrYkYhp48J31paHhCHbnvNmIY6vOiAC/AiQjRtD4l0OPUxos52fGC/6
XcnLldPHn7AadbMo/BkWIVRSAiSsw8Ta1w+ONb7uHPuksrx3DngE/iiVYZk4ju/jalS12DQEN86W
kHkks6Vqd3lg+F9uhKHZz1wg7T/uUJ033MoYn/PmroSZCcnQgot3fr59H9njEUBPtQSks7n+iRWF
GWP/owK3y7pS3uU8yx4kdcITft+lyC3Y19zBKrhiBtOqUufc2e/d6hxk1VTCnSDSTEgDFD3JiATD
7utHsYmn8ml7eK7+bFOn91310H+hHFpzdS4aVkZjqfgi46EWuEhzpEHfSDlXLQEsAqNJbB7ixaVK
HbEAVjHj2BMvnnVwrdwWVC72CvA7rfbQtbmxC2MIt1tKs3GoBcrlzmsM6GIhZFjJYbk9m6aCAbFm
oJQRTYOsgMH7S8f4X2VNQx1ssfw7u98W9R+YJpJtvEqXyPR9k57jt1K1eRabFpIyLKmfeJHCX+YW
QssaZhQs2xFnSXxHSlnIW9kMBLWj1jUwpqTjh0xy6lVjP1H4IRgXlzI0FZM2qMXsEBIMQoZQXsFh
6LfVls7sjESgN8+xbRGvTxZjOcYKOA6H3DjNHwtxsTMF5zOOgLsnsQNrXqpqqa6dgYNimRytm+2J
DVlFMNabhDqoyDDHkAeXFjGT7zjr+V5WXLSvfwzww9Yw1OTVreNEG5mlrz3R6fKQAASg3j0vdTBs
/3Yo/gTl0rzvj4oZnSmlKb7iyoyh8pGZ3H6KgXSmhzfanLbOmyMub1SKufA4vbR3yauSbUQ6rfss
Yo7q85aa26XyYguKrQ3p3CMLif91Py5HlH8JKru4EJnnfyrRZBdSR/ye2UuJWL05DUOdZ0q6HQhi
fnA4s1SryQNq2UsRJ8yeuW0pfFdIjX2xqUDfV6Ew6uHQaLSukV+j2K61vqg4fReCV89xENdSKzuP
3TWYSD4fMBQH8m9Qnu0j8iW0AXESetd9t8P1Ul258VgnFCHvU/ehbl3XRY6+C8vHnoBy3tJnqa3T
twQ+Ld/RTdnwJkePyy3yFAVX3enUBbkQFsAH45aQkNzvRtDcKGr3My8rf/Q4CrNfFHBXXh3/lAcW
n5Fz2R+k388H0KSfQ/3h/jUIiOyprMh5RscJaeux835XK/+6L+YJb+LJTWz9mFw4fOFff00Qv/0+
9wwwLkPxrE9nYnr9ptSB9/lc9euTqN6gcBD+UyBNzlrdKIe4yTup7ArjMHyUAZ2qm5KXCxI6qUu2
OvrvaHErVw5aNOB9VHkd4E5W1t0qMhfu0j60sRiG02kpCngcn5OLIURPYZyVdTdy6dO1SoX8ZCKs
ozS3b6RIsRBYgM8F+b4BoQ/B1lJEIdqegfrNuMBqQwp8E+ToWzltVwtZkoKNX+8l4tuYnfDTJ6SG
tpiivTshpuhMSj2hEYOiIaDMILUcmJ5sZeyZ8d8SbV364clMQTkGZrfPwprlcIQgsD9DgWiNpWdF
Zvt2d8Bv4t8aTWRMEqGAmYuTUrcigVS6fnJOPGv6V3NyMheYJRSAy1WjaSnxoYl/lRequRQZSuLE
Y+TJ5NzhkMtjIZL9uDv6Ez1iZClNyoWMuWBUv5USIiaUpJ1vtVQ/x0WqvIQuH3E/Dbo6CFS1RCB9
5ViPHh3KkwNmz2+if0PJJZS+Iyij+7NO5zLtXRZ5JmRXAXn0lGWQHckJK9psLOAy4jkEhq1yuflo
hC6+I7ZhOTd0NsVU3c7C7UgYeNYHmNoETksfBcesNK9aFd794yuKy+S8UwJjv7aYMqCFgXF4F840
UuHOc73zgusc75hgwgXqnowTIffoYMLlE86so/doH6MUZX68+EVfM0GrO09e61Vwe113j81VDuEK
XjDGmf8zkc4L5NeOTPdyvHgRDCyP2z2adn8a3oxHQgfJACLdeOJBxXpR0WA2posEtlY7zoYwCZd6
vpSTXjibb3rcfygyB/FDE0xHBUH/9t9N8gImkCoBa6s+aBbtLTm0gmgY2uIwyQ/XtoqWLguskk2w
B1YKhBo1MCPhB9IMLyGzRRZg1BoZn351goxWoFxtP2VLWnvtJx+0JipY4GVAignNNPGa1J6EORVg
isMWgoNDrUuCNDe7BgjdS00hNemW4ZQkqNG2uYgBMjHLE7amDiFBdhNjKTX2Bajo3lCFw58p7wHI
8v1nWSQLKJy7oIQg5lnoSOlwJDrkVli0cKIaYAFPFeEoN6QtIFniAWmtWw4DfOwJHq1QVKOFJeJt
4NMrHssebmW9PjJ7DuID2FO4mbZpVeKjgPW76a1I/8AFesHXNC7AvqBfaEwyumdK4Ziz7Pd4q/nD
J41Ai57rnLSjhVcHFekc8ohf/SbTtfbmQoDaF5yRR7QacgrfWlUwRY19kAu9+6RA1JOa2wGvDkC/
phCgmNNDhM1a81uxrF813FGuUhM6qW+FA/fPKFXKEyk5E9lP/q3bl2s3+5x0e+YmheShtlU3z2hJ
BkZWoZzs6yXENdAC3WuU1bM9CAmcx6Ie5kEvVz2yd3oqZVc2/cMCndByO+icHB5oYAVd3y5bbANN
MHSaqiHV7ANFMY104GZgcPNSfKR0UtPIUmoEuhScVEwIbyB4CoSkbjyfk1+tY+TuHTLc/USmiCCS
rxbIh+vCZuMqRDg4w5tk/A6XWOYHJgznnR6UsI4iBysMK6Np//I0tVarTto+/FvMa/WloxKpCtqj
ujTab+hVGILpqFXnNoiQ+8K4gDrLAr2cKOHvm37WcdG7p+3yjg6JrHVsRqFNNOYb5jjPXiJzMeou
YBgH9uufGq+yuijqvAsfdjVNtGw3ThGhjBsi/6o/NPj7oOUQStrhG2sGGT51hdOR2CF+B3skduxf
3XWIhYFQfhhHRu/kyMwgCb8wznhTb2KexOSVREu7vs/Jqm9im4dGncBhAJCTjBDWd7w6fESPexSJ
9FvzO5mYXBvNlWW7IJsyxmEq4PPgP/DtuNYi2knKpZUf8/3ig91RJEY1eWXom/b71lS1gz2lBilX
TSTvtsp7/FbXlX93vkVG8dOmiTGEzEX+9u3QRb5v5/KkvGEL5X4FtSRXnfjF33xFt9i8jvOBehnH
muD/ezbbgh1lAQuiqp3KNusMBrJ3doBHBCNorIFtqKgSKTpG+HrdUit/CY4mAsMHnQhUs0jSFn9k
pcsOmLtwnR2VIxfOBXjKY2+HU1W1NgPbrKsxWUMm0UQxFPGoiQScovGmVuJt73fgmo7TNn0P3U3g
TdGOLXPGXTDMNkpEvv1w9ezwml8cZQ/5BncOaqLCk4oWZeQ4WRo9JMbS/OBIA0nfuOFLGGfrPF4S
gW9Qau2gPINvh/wjB0G0RiCEs1SWn7hJM1uwMOjwFRe14WEbtM9KV/bkssHmWNYQPzjiJUt9m57C
clDCyy7ZLh3nwmZjONEuvQTkkaKlJWEa+oN+npOXbQAFDpeCSMCjpy7u3zjYV7i/kdzD+iLVII1F
Uqs1ug0uH1LnEIar6K6ZgegsXWV5CBog3kay/bXdyFK8j5e9hjTEgLGBSRJ9gdlAvuYs/M1CUJmZ
GxwsK0TngFSaDLxMaoRMD/Pv03K2JAgJQizJaHLyOrBzmBnXVM1C1ktbjGwptcdEPXVCPQWwW/qf
aJ9TENy6FiWoeRQz02mB8hY50AfCOeFcf3IxekzxnMQ37oYx6z9B9aMYqUz/ypIw95XjwLH5tS+F
feG8yBOorcn30B6//o6KY/cXL7VCf76H3LJTJdB7CzLPFktIsT2zE/yTR5wpo6kwyXGQrNpCOWvr
OGnRqQ81RndwGR7cJisYxD9Tb7gkGv/VxLNGPDaiBlpx4YiT8M/P623RX5SP0GWLukSCdwS2gmD+
gy57JOTMI73IEN5dTbOQrd41MoxsaSCN0BEFNAooz0mMV6Oqn5ZC0zK3qYe8lF9W+1UtTMQ3csxx
g5AfYWzP888Av5MrDwYeX8hQuG8igBb+t2M6k6OGQ0Eh0XqFez3/nus+ZgNRTNcvu3M3PouhrXmL
D+CawVEf9CEnp+Hb1G72jyXm+FiXIjAqedvakCaac6FIoA8NS39TV0xg/AKaOKp1pTr6c/XzThuG
2T8vxg8GQQI+jSnzRzL9X9rdOYTAmzcHfx2sMIWLEj3Ac7AhG/kzs2Ax+5EFReboTNEvBYbKtc/G
wuAqMqczYZaM8ey56UY/piQtWSyQ4BO85YPBqCmUxCEcN479WOnU0c9yBIB1yMsambIzlYH7mRTc
OmCb0atb7CH4LmvUYa1To9IOVbF7gQkiEXeshJgm9IjWpoVufWzdNG8IZF/wi3SdJYNz4Q6wkc6w
JIyr3OUUskuTrrQXyzFoDFrqq/EC2Cngkg/dAuU5GYL0gSs3GigVGR9wuUlNy5w8EilpC+ItOxEp
As+/ulgPlLXKKaaDo/tkt9Y8qyoh5QQ/RCbi+YsG6bkrvC019aRsKOwqaw/KanMgOne4i5krzoRF
Ke6mLNxho2JQYFn7tCB3MnQ2p7cBziWQ4l3DstzhI3ZZWgZyywAdxCwYn4j621IwbxwfyRMHEi9A
BexJm3ltI0FUzsvCg1oTJI9hcGW0I5IaohcY69kIZQzH2xT4cRDfTJ84gsyitGMcR8LYOI5CQYqu
TMnDoNj2770pgCwtIidl/67reUL9JPmh6zzHzPCXEJAGcDP5CHKJrQdUYlWb2wxl9NC7aCKUABKZ
rfuWQwvgahJ8TJr9noUkGXSpbEGeySp9zaGRO9LQ/bP78iD4IhPI6v59kVIYFGSC5geJlKRy95gD
y1Zgi8+l3wdUVALcEEX5lD2CIu/pyC/oBQG5IZJowReWVHRIAD3JfpqCi75M+C8h9bCgE+UPSaKG
/U03r1yZxgouNA952fhDr2bIOMaKWQYqZFEAazoffP/ZcWZXOTXHuwKzycPEyjlKVXLS7jx9a5jb
ZajicyWZmwSZJFMarEJvCusxXMFdb2TlDm30U3S0lZWB3X74sbmFecp+UoffkuPGQQy36eZDGTq4
5WH+G1A3C+sRBc+r9rmbi0kCzcMqR5lquhOjxoUX6FNUZs884RqZpEsPyp2DLUH+OTNzwA/Piflr
eOyaL5NUZFavLo1yy+Cb0FfLUktywUHRB1LdvmCbGuzRne9sek3KZ/VUutQQkSuBOUDTL4h8qlDG
7YWgqqugxdQEKXnkabvn+5xLUAKuWgmCcxSo8SiRaGqHpfVGY/ElBl2Ixkn36P2IVE1KUPDmLh3V
kqXQTRaYutbaN+HBiACKX0yMWBRTvR+KnfDrw4ZP5Kk7cQ4jxohLI27J5bFOXkoPwgoTkzY33ILk
FzBfuhVSK4gocfMZnxwnUE+1oXRy74QIuTfZ+YqoC2x38rEBIR3Ffh/cuEcRwNR8YRtYMP10JVct
FkFq7/Th/VZM8rYROQ1RmdrUFDbJnF2fHeVGPt5ISsk42wGtvTLGsBjH1C9aI6t2MDg5IFXjuWDM
2Q2aSk7j8Xcm4obowFbwSte+cprcOYR87cRZ7v1IHvcYCnA8ceR9OlaLLlNPRlaF9wjVMATyIKOy
2ypM6rhf18aLX7MSmh+qMLiFL5FKIbGQYTvk4UH+N0Wct5oVR583JBs0QGJOF96KdGDACkQSVzr4
2QWsUqNpw+oTE8SXW+d+F4Q/HihesPefU7gtq/3N0llz6iaz/IlzT2hT7ow1E8ZjvfF5EDWNLh2G
Yy+Or0kI8ZSi9vdPm6BJ+CEsx12Tvj085SjHUoYGm3z4HsHpFUHN3qUqvmX6JMC8aQMyWk9jdZPz
PDTOzo2GhCwjPLuhmOAHZ+byVFSA65cuWGmrs8Arazy6dR4qfwvGteEvpA9HIcJbMEffdTugFtXY
f5VDUQN3btxKF2frGzmDHohykixCUveGLW48YrSJklJ3DQsN9Dq+mGr0HCq3GNSNYR4xVs9kMS/4
EKoIsdaItbrQHtO1mPgYMX0aB+aLRP/GJd7YsIBpGvv0zqdq8BrM3VLdl/NaxUAzAuJGjOcjP+ql
aO1+tHi4e6MB1mYn/Qtuuqr0OioeRclrXc8Zu0kpfhFqqZ6RqT5EQxDg55xKprwOHUCamXiW5pKz
R7yTasgMAE8H2F1epI2MndZagn/cLTF+XVMlBKFFMcs4hBqDdqNv3RpjYSacRGz5Kj0CCDxbjrGj
LgliFqlmSjLvq+pN9tm+8SMKX/PMZ8pW6B1Git2oZJzmp6pHYtcZSx88S8M5N0GBmidVcJelKlLM
wgNzI2jqBIW7zT9WQ5h9W1QWTXpHzbQuQCqMSgC/n9kRmmFiHHB8LBJ2+qYTkpBa0FC7J90Px0CQ
weF4SBfuU/cWQiYmkD9Z1JYiiWXLvVQq98SBLQC+UOS2Xgroa/eVHPH8dUtD34CnHTt6idPgygBx
yYlzCVPtuRV5lnASDUhta7/RcPQ3OownnaDeGyrnq8RaNMHiH8zfpz5Qc/Tk1OYo7wI+T62h+Yya
pf5Qv4q5dINj0bqtYIlpq2O16yoZ8qJJ1JLQJJNxjTTCcUSfXRMcfp2I8C4xcl63Rm7U18kst+SL
i/hq65dv6s1W2ZLEmNICc/iPbq3dsZxHaZ4CFWGeFgJQDlNAEcidVQg8RdQdeV8RXpyzxRT3D8bo
MzdGfr95pITv0TAueX22iXTtfEz5IZILNi10iZvkBpMg66swydo/dc7s35FdP2xek4joZzhkrG18
Egq0t09veGgBptXhDcapU3qeoXeCee1A9vFh90agaNLCv2Q5G+TnX/mpvjuiFr7FS43/JNNl7MYk
AaPhAMhW+lNre3oymT3KGauqJ5zhB8AKACXSUdx3hHqIaYXGmWp4mL/SPS0+HwXUhW+sHJ7xVrr5
UIJBcZHveEWZbBuImoxtN854VJxLfJe7GOZwfBWy3lxXKSXsizcgbFfjtD6+RgtvFk80pYFgeZpV
X9iwr1i0An/rwKJa8oSp5r9aCoMca1zpkbZn+fPijL9+x42cE3oW2gl9HmCNVIrOrfq8nrgJU8Lu
YbbMAp0jFWxsrawJwIv9kji6owt36CL5GOK9wc60XnWbqDDfJDlq9lXN4fus0qExYpRNdZesew2L
xI7VPRtr13ixB2jx/nVfTDuW0/HSwIWVPn55lWZup5t+wOurgphhC7IH5ki8Gw9USKXYJqj85yI1
e4VuJO3nGp0fxE4AmQeaP5N/Mp0ABI/rSVZoyT2Y+mvpgYlYRg7YoPpjJ3saqsd7JzvSDUEHSYC+
5AnfdFJfpuF9AedbhEWgPTpDtf4QwPeev6mzjn/hvjnayOdpPGmD4cF7bzt1GYO9LKMFFyetTS/R
AVRQl9iHAQAVgCUgBYkxD3bja05TIfTpR/rgfiRSiOfk0mmAT2z5p4SYhvazCLpaRz+/oO1kIHak
k+XUVrKnXkUlpXA+Z4doicHOGy8ghh3GqYMe5EJMLz0qTxjCoQIhD/OE6oXZgAQcoXUYtotVvCp1
iJuu61aYLatmIx06vvMAf0F1E2W48QATgsPPxgvl7J3obNnnTM5ealTFl3YeKMvxIqV8RWxyKNRR
svJ1fnPSjm2enwhCg7nvFIhMNe6juojpSJH5B+HrPXhlRg/WnWptyEdFuJlmS2v6BgQr3EyLuJw5
fmrxM0a0TJSXOgPSrmHDVwGeuKup1tmyEIpxj193OdLGOeyWsmPFQvEqNW+nboq6QicZeKCMS8Gm
gSKk1O5apMELzuXEnJa4RpoejK54mpbg+n2dbzBpWWuOic9+9PgzAa74es8es5lZ/T7Op8S4rTnN
leLtF8WXX7XjlY0muJxCHtMhivMmKVLtnbzPzMLTrca0o1OF4cHJuZJjSYM2sDk5c8qiSSHjbnKg
uKiYY3KhDVLpO/eJMTqg0DZYUdMwv1o9HI3sOVstJUEz7JYuvmnLzovug282YVxkiYISxDJnXrHi
xVRSQotkcrEsUa6cSY2sTvP+orW1Xa/QkLm9DDm0l/vScGAxEPw8bItS3BHqNPkChloEGzT5pII7
WUpnsNgAlnNDVTP5SvrbfrAAYjIv/E7EBDWzxJ8US30hwIAd9c0nEDHdV5iDaeuEcVzuKi/z3ykF
FXb/OuG/CaRj3zduoBd79fNyQZNFftW1B4uwdeOq5cmN0QhvlLFVD5/cGVb0LyAexrAa8a3P0vsF
FUUIcjPwUUoAghTofFf4mZVFy61yM3n11+8EkRuuD8ufPDkLIhFd9T0aiTln2pCCDmUhMnV1z2a7
IV2FOP35DXKmQLgGFmFDeSzkV6IX+UtG2H9dUBAMSCD0zDkDHEBDPfnRa3th9IvnxaO9joTgsnDo
VwNveKng0dZydlgXDFmRAECSuMnjZKSLWe23WtG7Y9l7NZyY1vYTBiOJmNYPPi2BQRk6fZ2WCpCY
qaRzzvzstbQPa/sl6BJAI1wqe/Yh1d7d6i6gZRp7XzznT09v2KS7sFJz4Niv2B2ZLJAqE/lTS2KP
4tBTUx/lNeaY5fz1KEfR6QhCngTx9uINkobKvBuJEPAhuNNe5SwnDN/DwCeovTqmMkIAs6ZsTKA6
Kmy6DLx7vSvH1F8zqnOAuffXwc2gpozpShGzhlZyPBEtXAfbhEQEjiQ02fyTRahHkZOKc1VJ0+56
AHyTvQ+1MAcO/vEBNnh1CG4Xyp5j0PWvGWwkBngafu25tE5T1OyQzTfrMj00RFjBnF85AVLrVhYm
6jrMQ51sQiHVaOAMjwDbPbsw35D78s2hIkIJiPNl0G2j/w75rau39g+5XXGSRts5z8EWuJXTxpdF
xi1tWfPMI5keo07S8RE+DIgYUsUSPUAy3ownBAy6NaEYwpDA8Cn3Yz7/XgoCDK7qUwwhUQ7ZOqqw
lCG+LKo0GiMOcpzbZQ4PgroQq+8aOmQIldgEyGT6gJtI6qLn5t7LOnIqBEDN59JhvEiQW9zdPL7w
WajVzGzEBxElJeqgMI2DicblGtKNa0BadZgfILFebmoHVbzjv8MjCZLbuuiSJI8sq74At/iVcGwk
UhuDNcJ6Tu4VHcZ1jcRV3lrGB/YjIXRMJOVnG+cA8nfmrGhm4wbNAKTZCIX9MAVaw3Uskruz4K67
whEij2b3fXHLUxxJTpKhrYC0DhIQhMOa0r6PsZTapX1NAQlaSAx1tdp67piPjTOGlIamn4iTZMTU
nQDRHaujlWtnT78UsVhQ1wrkU0qQbLi8ZihdMqDnB+Zcq+8L5kWVXbjf/Wg4JHbSKt+jVSwlzDs9
eCOwV3ZE64faziuosap+1K1JzytX1Y2X/IFt4DHY6JokMRKVGQ85yamODEDgY/qKIVI9dR6OJanI
+Y6r2/YeCec7C64UXyyj9Jld7UaBpoHTHuP1E5h0gDC3pLYYP7gR79ysMgDn5ycb1bi/9Mfa16LJ
ovmX+ZaSgMJ0JUqdJrX6D4S4pb7yTjbt8Bc3R4G+etNdF8Vz0QWJX3z+KCjcNaTi7TgjQdqVj39W
mwQTWqAM6n6PEyFO0VlnsId2KsTqRsDpMo/oUQPI8psselgKPy0+zJ3PPVYRIXnAghJtuQmOyTOI
Y3ZZJ7FTaKra58E24QfFA0Y0hEet7IIphaqxWtZGC+lMKOzk4Ms5Ymlz4+4AZcwchr17hs+f3XIf
eCG0jorjJ+fRlcHc2n9N2S+FIGPNh5yPBNUihzkH+v4ykVgYlJvrl3SoS559GGpUDVyHR6vCAd75
G1S5m7V15Zms+tg6ky6pM5lK7kBmtuYWN9LEGyGMoJEArvL8NImxqGbaVA4AEsQJbSVeKhyEIp1K
CkcEg5RE0ZFoviZvDe3B+oRWiUWsaBe7xZr9iwSFuR5TQDRdNOpgzqm1czLkapCdYxUncckhY3qN
fY8yvNVNnL+mxKi4J8qolQwaTSxFPRy5jkEQvSvMuzoipFTdg0/17Spindyi4LwssIJYdVgRMEyq
So+TO9yZFdanfCaWUZPFG8RUeZZdYy/tG3QiPZQXZ0dyBrXRT/7bFiViN6Fp43KaNUWS1d9IEsoT
/PtCE8JElxbCbRcAIS3Dk1li5vgI39e2t2oEesspvAAc9N26h1HGD9L7tm3RlamN5BI0sAEy7uLZ
UkV+xQMvERBLm8/SWSzEMRnln+e2M6z1cGngF9Tys++L8DNviWeESaZPqI5JHjqpamulxEQlV9/S
5SVgtMffoJX6Yb41I3X1/tLC0jNITPGLiifLOaugUVmdKE+BD3gnY0Sl1LZQ9lKNEKyVhL3OjmN7
h0pDDz4G+kGsH9v0mU/434aPoenmoDY0i0PcIY3Jy4mF/Hi6/JvrNt87lKptR6ZA8H54zwmsXFzw
DHxMXoqbPyNAl8oFos9UjWM+CyT79bwRdu+Z4wLm0nsGRBtQsERu9FetYbU2QClnary3E5ObOSjS
aIyX0la715yS5PlAClP0CC+cpDKsHUhsMbVzdzH3AlAXCTvufuoByjXrKcyqnrGAc7gbQ9SBx5Ng
QFLibKMeY2DszhK7diXn8OAzAHeOmR4+jnF9XmGFSXuXk1F8KT+LODnnux2DUWZRT6xTcBgGMDE3
bxqtJySyTwzJY0FdlCOTXOfGYLJvoshhyCl/xkEjmL+KKfjBUsxjKLDZx00HZ8uwYzqXckjSCxEC
XXE0NfvPtIfO6EBu/LpJEjtgsHEYG/S/V4vDuyPBzdlgmKi96JZaQ/8p4iXPPdYAwHbapOH5YKlz
vHXZtsQlp2IPAW6WXw8Nj0YQhn4NO42rAOoIZwuLdxkMev4Pyv0gvSxPg5e7HPRw2pXGbVPOxgVf
00CK3IujjdpRy6nMMAG0i5NEZJRzLXgWf4xwqdFJKda/UxLyXXK6+zvY41hbl8dTKKF/NkPpK5i8
HpEMiAWEV8WhrvThySsKr8/E/P2nQ9rLsLhV+/+J7NAPa0yqoYoaY9O3fltYbXI8MMpJJdItTxWH
ghd7BoXS7DEg/gevxefYekSWT9UHXGQuSUTwiM6bvWCjwccDZ5+Uh6slyQS4cVdNp186P/owC/Cw
I0sKyyzrxDkU3J2hWh08MHSP2/uXE87gSQAhU1mjTxXWVfTuUhL0BvQO/+3aP6SC0btxL0+ovLZ1
efniwe5yQFJ0CLI++68dplh9fZuvsajvhewCAg0Du728dv4FtPIWSxZzMZacdpPffjtbKzAHUsc0
wckFbox5KwXeeKqiLksIZE4XiaGr0B46Z0HfpqRlZCbbKpTnsz78XKNRRlGExTGsUX8JmAvH/axp
ANE3r7QnFOtZ3nx3ARJL0lbKWrPyowvXchGG4z66BHAgiCdAccIawAVJArlLLBkVOn5gdmfOHCOp
IAOSuIm/ZYK2UGm8S//31itp9+1qFoQXiXP//bVsxRrisa4JYwVaA4ND+6uele1Vtd2/SHwY0Kft
+vN1zdaXeWosOXmD4q+PEc0fmL/MKT6BeVYTZIc2+/AG5AA4lFf3iim1N2eH2He829yeEKLmGMjL
BaiLO7e1AQ7YbrAvymm6utx9rPf8/Sk5Im+EyidseA4dIc1g9PUFqq2v/iZoufaxtLLdpsh0GAxA
VFlydgPdgJGNlm3zPBqfEPF15hWWlUkIkS706YdR/055/q06buwB0xjxCZmHO/dyCnxaU9e9xDY5
u7Ws151d+auHhAUYqOjI8CnVDVRg/q7lpf4tYKU+K/qW0eGdxFhvyzKIdnjBm7+q0WRxhBMGO5Bp
z0U6jrYircVAw5ao344q6lKYVEyRgB2b+tYpybUIY6tfqHcl30CqFndx83Tl4zXX1RFMiiRy7D2g
EshZM0EkY2sJU+YeXG/xal5Dd82xiKzrs0t1eqPt0GSmL6FfWPbwsqV4bw5u4qPqXkUqL/xACEPS
kWUjpa8Mhh6YTmYQm30iO19K9dOJY2yUYZ1QexPnKOo0GYzQZovxgC7S6oBIp+4lqWQ8vLg3/842
A/UXzFidO4TaTYLDOC5eKCYmIS20V1sN52pIe4mLlsYiI5alKNdzrEpeFtomIc9+9gjHfso2PcmR
NLhw38vf1whTi51PpWQN0h9W37iAcRMTIpPslaqBZrcWx8BYlai8/OX2YvLiT2wHkgJTefqv4KSL
1PcMy5qw/FbcwSkhRoaEyhnFCL0PDHXLYWOga6mlZ8JS+SC/0BzrPPem4iDMIQY3Ie8aX8pkV1sj
e0rf9qkf1+Og8dTberPyFWeXPN/QCdi/oHU4Gs3/8ISU6MWrkSVju+vGqtTEdG0KPfdE4bjZ0Z9B
4oBTsKPTO+gPUC2UwgKEx1eifnnMypu+Bd6y7xJsAk1WUkUEHQbAy9KgvlP3UhaByX3ANI7/B5Km
MMkEHjsygQvgQgArU1Qaoyl/d7HmM/cqLIylz04Sy1ljcGTaxQkX3O5U6GCOWMiO3GgS6BSd0Ywh
99clgL5oJYWgyMtzC2i33kfLzqVdZhRqBGycNjwK9lIshOrDVFNCVZ+msumJgHA9UJ5wPHDh1+I5
WV4Mz5oGBuKmNTWgBUtI41gqrDXXK/xV/iTNnubY2RDIdw39DdXXZeHMu0szA4CQXZxAjII5OJ6O
lSw4fTBRFB+OOca1lB7OPmY/l9EwBrNEWQsPluan42hZvfHKJKx2jNvzRioRZrtwoVsNzcfp2Vl5
IC0yMR/ICqjZYxHY3d85GrZIXH/d+XXvR1ISkcp7mMv1Ur5AzYCfEzKPp5J6FL8XuWhW9OFopfaV
bySi1FT2xKijdKOITrBJ6fbWqR5Ics8zqpnnzXiWxcYGg91lzF+6us+7Bx4c4p06nAXMyHnmjaCc
MWMe5hY2VVxeEDeaCcnsWC3WEUnqut4w+JxAELLidiTj1ah3xslh6NDJl1bTitxEx2DOryHln0Rt
qfG13W+Mhwy2vVtJoqYzN47q2IiTZVqJwojV6zZga0IbS/f9sp3VD6ZJwxYuDhVq6rTUWnffFof2
oM3YzX5wHAUvr3AkLcHRbSpC3KIlQ/4SnbP2SPuDMiyIAIOAQi5WudUnPfpi/WkEW5unRhEwzolE
aoE34setou06DZyVHM/GoVijQgJ7kgyhwuNUfxsMuVgCsTdKEjBPMZJDIZJfsH9/NAYWJrejEEIp
VDobSRQ3w4puULhUfa/IMYSJ3rq0eaegkiayqxKtY/9bkI2JBLBSYeVTtOzSTf+rbLaDsZfjox7n
DUOXO1b+Gelxx1pEq/GsF3WH/eIHEZekKq0gXCx2gZF1hPVHwru2Izh/VW3k43AfggDcVieroqrz
S+VlZNJHiWcJ6xKAaKLfJF1ABBOB0QoKKMp3feu3aoziGbpdytdW4zO+as29FFEaigYdqwbC6km7
qQ7Nmm3zgkzBuxQqOjtpQu1au/R89x65r9tLgP/LDz7Oz3Y1uCAt0Wkc+WjCV+S1fs+sz0Po0fa5
bFq9bC/NowFd2TkxeRsuEMIc00OefP7QB2NrAXxTRIjSfYPBcp7mNAepsbWkcMWLnIsmzFmxCgcH
MufTuJVF+PKuIvNS4KyxS3/J3iJVVLzvLiRkwJ0RuPRiSrZlh2dyvYCM67eOA1RFAq9i9DF+IcaN
Hw5PB00BpEVl5qkYQ8TtuVdWgrCv7XaelLLlcDf4jjBZnvu0/aYDQTCXbwNvTS+H0ilfHXhYa5JW
bHngK+oWhJGQhc8798QuZbPShhGrv84ILXnfo53WO+ggcDhixmweS5dbfvD67zvthEzD2diTd2zT
OtIviD05lraCzOTJLObGQvYF6JSIh5x7KdU10imlSE/g4Jd0F+0wodYhHqOoajzulgrz2RTQEO9o
tqT1lMysWewOdBAo1FKh8G5v0rBXNxPPWetxuXOJu/+zAvFACcXQ8bHT/IMu9hqbRLYZOr+GKGnQ
AABAZDDXFk9LJNCTjza7BfT8isubD/iCYhLsgUii2wZcHE5fcFYJIIX1t0satoy9k2BtboSQDHrq
lbeKLty8JECtvbanyFbcoK8eMSDHKgV+2+/lNoeo8YMjf3NVr6CEWK/Jt/0rwj0mxpE3yX5uU5xE
49zUgJdpHxsgUoFzVyUmdSFPTjqHsdFHRbSxQk/M+fRUldHIVOImaPCQ+wzoVZji5MH//WPRsPF1
FzlTpvuQdBGoF3t9oG8lZF+Txspwh97Z+GnhmebXE2GNNE3yA0A9B2LS4xap676YtlorzFQUzDQz
RTDci6OoXeWk1AmRa1vqGMiZPU9pcUwxx/nHur1I1zu46wm+ajeDMlij92/HVhHy1QA03UULGHYA
Kx/5sJHYe2chrrvhe9DC+JtCPGp3pMqIoaa8JIVPyzAZpuW+Zts5nBu08AKIA72d7CNPaYkBYeWE
3F9B1BM8Um0xKdR7HuZd3ab9iwsTbkojm/vzN1eXA7gVRYqx3KN8kAlUQkVmit4W3+s9dD5k/EU4
lRVhdSEKY+2+QINRF2WABCiZhvMufM9f7dfrEXnJ2KpFMF/s6De91UVFFadrJbPPe3ofJZZL6Ly/
5veeTqPxgnrK4ScIknu7d35itbgO08+QLUM3Bud+5PkxWGjILb5V8IomnHNPSqdqorc/rRSA+4hc
FZSxlNzIXK7JS7PkVT1HCidxLhPZtK/1t/fKhx20Xvc03UHDx/dPNoquyJONoMIxXpKVUsY03/e5
OJT0LxiWdXCC1mCsZv9+4rXi9t8upPXFU3VfUy1lR7u3VmPbFINy7k4QSVH+Z7dr7W7Zscyqizx3
n0v5GhdiYvPOXOMlCm1arGIowUX3FtRrB7kq44PzfOSEKDPeyVDbUMXLGG48MBZBeTHTPmI7R0Zp
wxCUKQIPZD97u4MoATv8KB6QHddIZzeP6G8o60tCrB2DbX+BsmHFsPz3dkiDv4bN0mR8msQAwn+K
7MGlFDGQqoBUS3hB7d77m5fjaDBh2cu5B2cwZXFUm3F0ws897ZYjdDWMfw0cb1zUJo04sqKKYuHD
GavjaK2td4RRr2i59tOusEujvf1/kNlp0gPfUZnSUpAefwSk+1T0PMQHrEs3PZWWvny9H9WjsVea
2R2tRnNUYRFEN7rlXb8iVy3CHLmd0zIUrRFL5UNR0sg44OXkmkThYdfWT9TfSjMTa5nJaJPfI9n1
OQOnK53q5Czjv5vsjvWPgob+8y2l8ISEVwSykoY5zmxMsb0VnfPKTv1nyKThQmzfztbR2s7GbJOR
BKZ26GVdqO2Q6U8foC0WyPX95KxGLzU/f/03g+aohLC9JoKm0tvih28NBoPSVUSPtNKLGxmTwJTs
nzhE2DVuJ7d/BEQcDKAW1lHtior0W4EUqfSUhpfVsQsbrqfM9hQJc8zkqYHv63ikIwgdcw0wfEFe
k2G/YXepTJpdAcLhccis7yBshiuy+6MM7ZxxJ61LOgPtXqusf6vPGfcpDAM7YKjBUcJcqaxhHO3M
Ye0yBO22m+DL4m+ORM71sh7fOe/ScjGMoMIWAL2ymiTxVIDpz5FwhsR4/orhVoUopro16NIWLozD
fkuk9BCHYYLsvn4HzE+QxVdotMeEJyZkDEQZ30wGduEMiqWBrRIctptqiessxq/HDg77SXAS0ILT
G1+uR0sKlbQX5X5VWLKo4ughgH6zQLtC8M8kVM+U7ZvC4VKxJEh9YH+OAY10U2hmjdPjMMA8HPxA
I9i0xAa1ecuDwY5gpe2/ncLbzQnfYKuk65Xh974uW6ubwwRQyJi/aVLQTXpeoj2IPfdb56dL+UU3
qppSgmmhmW34tyM2sijuIW5eemLjqm1ws0YAeVtYpfQmKaLGBfQbkgNsvCWsl09lcPmniRf0+Xvk
Ke9GPQVWB3NEQp3MOocJMlCLB/tamQxlLOLFC1NFqdNoE1vt51OWJfOqJEiZGvxgKd7ZUTMwtzWf
VQPQI0p5EtYEQXrlyER/Mx7uXdZm9wVzhdrLKB1RPdcoubSemaf1YVUsF2ZY3ObwGOoecCCifjE+
RiW07faZphZbiurn81wVOsTL2tE1jhDTTzU3/vfTxpcpykd+d9SGJqB1WKuNfOrghMNMq35KYdWO
38d4gtICwnsfOlDz1eQ/3Qon8mpBGPD8qlCOQ7Xuo1yJj228z6Kg9Sw/Ec7NavwSpSN+HXgp5WbX
Pt6zi/fwvy0HNGX8GDVMQlD94gc8DcIAHrcII910IrKnBtrL5O0sjTVJG/rDWOqi5m9mbmmlaQdv
N01fwjt4Reo7DaJMUR/z+0B+HxlPpXS+lUHWjkFb+0TLymKkifVLY2Zhvap5Y6Mz0I1kAu682T9R
mzij0AE2svLRnFZJVlKvqWAYOy93i+D6vfsH/pZPMtwSasvpDnTF7l2UQNoZSwzRBbcsq+HYQWDy
i8txC9oZEX3w5glRMifCjJvA3TUobb7iqgzB7zjVboSUjksIEleu1Js0JSQ4OVNwnfup3GHeR1GA
XHWTrgzgbi+9YLEPLMfaiwTJU8Gy7IBWkO4gXNCw5jZM7/jGI2b9qb0IL1wUN5TDfvKh58wW7DUa
Dho1sjMAyFUYHG6sP6Tqq7UASBrBJqTEHlGBWOm2Xso74heKhwaHwDvJIqMqTMr5vIegXYgELuD6
kZWE86T56ebs190ub479mG8g2ov780OIpEfY/Z/mwF98P3V8bYeDgqyUHvAAupXVPA3cRnnvnSfd
v5sfNbZ/wxlts3v4MjSIM+WJ5E4BU1JEqyFTycKrFXwfnSmXK9iQGCKFFPwp9sYn/RhkPIIggw9R
OZHc+KpzSni/8LdUOuGEr9UyWn9t+beTpVt29TYSAeVq1Ub+PS4QleMl9H+8fJBZ0cdWZvVNTD22
L8/6+sMD+HzT4H9fdoRorKR4qD55aI0OQSDg4YISJAHxx94JJ0bWypa5hd9Z9h3joSLdooAmnQJj
eK6ZvXqaGzySLpRoPIGXchNRxpuvVnyVjeeMPcdGJGFxY/kvqj+1UbttjKkv6CKAxkAJ43hmWZgy
1U4MD2pChPc5PVwuF1MkJTubYPf4BHX41xKMGipZC7vUrIvW1jW6+UqfXBnW6sGEtVbV7d2tKaly
gsYds0/i36Uascb2iC7IFQP39J3vhwjYzbayy9eS/cWvVjPAYiltoMMEjee9ToFT9XvguKyYE33u
ouaNe+xNlUrVSzT0uu7cM/srdNzUm376i3tbWurkpLb3iKyNXEoHvYst8y+dBhiPzChIDokmFg00
VQW6rst6zq+LmvObB6G5KUDuSFb6QKoSpNNLzEGE/B4gQxKVBs4QUDqJHlKtJx8sj8CRofVMYXXq
pkABKsDP2jCr46zapAC1M53006ZtU2/vioJBaPXb2RrvOlBA2gNi2aRkzUws1XSRPcJvr7sC7H3V
jKalR8TXwHJpGU8TFRl7enCX4L/Q9LZjHivY7fuWc9tN328dU5hJ/slGilgpVBcIj5IAwX7Bdqsa
mFriJlBEPZMx6J1qmE9zIjJeyoEWFssNFJ5IMBwVQEZwnNLMqoLCQv1ezzFT404J0meSfxdh4Bv3
1CDchVHcyVtG5rvKmpr/KyUzKY5+dtw30YSVBQkRtmE0gjkNjUlXW2P1W4j/M9AhEMpB5tm5i0CU
xRCZE9xqTb4oNgUyr78YubMXyNKbYfGdm9QFzpvcXG6GRToRzgf85H9yGkAzIP0Y6n2xtQTNV1fS
L09wFrk9oJ3I0JRm8uezvmgFbmL8ID2s9HK6ZYsW1NxTweyUjYBEl0Zzb3FCQQRy1zG0VS7zDFU4
tcjcMenlbmKIPShe7Umebkl7nrQQiwmIr/L+jTdSVX7bU8w5u57V0y2OI5EZCVyFozGwei+8Dp2r
40Nv4ihgAluLhTjufd5kKTUvzomfQGZM6m9Rg8oDhSzCjIIEEHnfgysm1XascCOkeTvYLVlyXAR1
Fl8700m4rufM7Sr5iSSxscGx/Hen03n/EtFxV3vejaHHsnmYeU6nmUcG/mmzTfcyc2wO5/gy3JBz
XeiOrg6ILfncTeufPTAPE27R0gKHot7B5/VnpOtUfHuixY0d3N1JCnsgoloAtJmhPU3ifFBSVNLl
lPR7PFVcMRzI7+FUd2Z50U+EbxN1Wb2Tozj5ihVstv3n+TXcSiVhMtcdAeXgx4jevKMNRJrUzdbN
uWrudGeUjPRXstloUt0lQPzSNj3u1gxTjTbPUkHrYve+oBXM6dQXb8w8MBXxAoViUsoXkphQkbCD
jDoGCejQUCi9a9cZMERHiAcEqUjpt7be5WkiVa7JDksMFfHkJrnAKNhohASH6nBWn8r5JZyTNgOH
1MH80VauDRj4rPNUvrZrbzfPZfiF6ZInHyckAhu7tXZIPxPFnd9KM/AYN9FI+kEG6gA6e1W2HgKS
WZqV3uFgnECmqx8J5NwhiBsH6Y7cyG0d6p3OR/2brxgiKpDuapLWztmjz0sIM6hQOSBdcVxKlsx5
hHIdIklC0MhN5O1m5fKzGYuGZlUqLYoE+Ny2B0EtABRmBQ3JN9O8KpNFo3Uf7+Qpfnz/2+SZJ2CU
B6EQwy3tBpsQ+9pZ8cko0+nx6VTqyq9Wo9tttSb6xvEdo+IYoAfJyDxTYzjWHJE9MifH+x3VB6Cf
0iuUhxWxgrN6116JfeDd2fQGt7YgE2JKdmOXZNNml92cplqcfjJncs+o2zOVQrr2Adi+xUUt1CPB
3EKlT+1L0fJ1BbzN37dDAAmxYWPLB+4ak+BuE/bBocNx9asYMZP+lD45akx77nal19bWZsCZQwyf
LD6dSc8KNrpokobeU/7ER08Hw41d7yZk3Mx+KPJZuaKMwgmh6dD4xCHyE0/XYDJ9lb/kX4H5RCzn
kFkyAC/ZULml5Dw+eO9bBQQShwMilp+xVy0pxx8WRXOQMLt6Aes/LxZoAjl6UD357wwfIbGq02Bh
veM3RqGDuP8JVO2EIYjhxWZqj47WCpvsu7Zfd89sKt7iFlfeTnX2IR5RwrRh59cA8ErO7wg3IOGm
1Cky9S4z/JCqVoRIuABQR13Kqxt6YPCTeUXod63LeKYqRVd6cFF6sFZz15aS6HupNYxZ/IbhYEFg
1PwMoHBzly6ltrn5/Hfz3kKfkdTuqgpCIw4khinzUUVpb/nLDJVPiGbam7fZzPvSae6+qS1k7pIa
3EY9beObQFMcNe8HPMnBeR3fizzrUosYe4O3TmyuzpWA7brQ9kq8iNDwqhHV+7Y82W2zCZsacdMv
dwypdiUhgJ06IQ2MqR38UZb6RDgCzb4X9aBiBRb0hhj8EfZOVWTLtu/WmEgPZO3Yeot5TEVhGQGT
5y99N1DSXSamot50qNd2tl0D8/pzoM7zYPq01+3onQZQabgvI5Zq9O03A6ZBUGS1J2vizc3Kl8Mw
KNod4N6HjNfAaj/yDo2tmI5nXQxmcU20aqACAFM97TjY8K2MoSoi5GY4yi5TjCYMGYfhBzVTgh3Z
TpUuZ2SSaH0aGbAD2a2soWQkxX2F8pfrW1yskNKJDmLRTC3P/bf3ScJhAFXtXVGKrshbtoedjUsi
pn7+AFGedTAMhQGmUobWGDyr71LRIoL1pwB2MBo6vAyb8K5H6c6pUVglaXWTq2/uDCgR8ioFC4wo
0uRnPt77BKVxANlQRs6YrTAWBBIcfjoDVgY3PHJfo1tg2MIivBcuf2Tn+bZAa2Vmao49ctKdkCLD
ZhYa8bz7XdhUmok1wQgJr/Uw7cfH/3MO8rSlPhhfXDkhtwuVzvi9/Mtfrqu6VISwl+91AzHKG9l7
H5kD8tdymM1u2ubvkDM2i2Nqwsu6ObKkKHJILenqjo2dmgROzNdPf/s2YDdpkFWD56+bfwZEa6sa
xO7g0ZRtzc1+g8WG/0pn8tTYL8+6OsZXuBZyn009KRHVK4qfDF/mRZKXc2LXe+aavNofGv2Q2+Wz
a6hhua54aSdFI77klmHZ/5IL8g6jcHoUQNL8lCItx90c42WMTjRPE9gbmZHH8f/N0OcrupWlJTFP
8FJdD7+vtYu7kSWGaHLNAEgUM5biLGnv1gYeVPnkZJ7E8HQsyHXg1b1gPT5tgEqJI7hI5zINqmwd
QyfpTD84x5Ubar8xHOpgMsmtjV+PZ3UYUKKbKkq9chuuR6DnY8mw34RuFIT6MSvPz17SumphBJv2
7Qfx3QpjcYSnOGMSvCtJgbV0/h0nfc+Bgil76fhmABtsief9PEb8ov6PqXzCdBungNt7ryHfh4Ge
eyNbdJkEIZIJvO9Jvg6tk1hBU9oB35cvHpXY4qYWrRu1zMc5tYyLQ4k+Zsmmr4njYD8KLg3QrcA/
zdpfAgCC1a3fpbPmjqZ6tKI0hX2+TmHwYaHBwkBbaj8v59wSrsFdPoCjj9HBIg/KW0qwZddjf4DQ
c3ssP+8LBVV/21jkPpQP4qwqZLNtxax8Fuio/pXC+LgZeTFyoqgic37SrFStNq2bK28r+lrHJmAl
PcIPOD/ueT0D9LU3ynsOPB33U6S2oVvGiO4KWdzL1dBQ/jz5MqWeTMgrvwgEW3vNzMDiT1BrvUP+
jiILkyZHm5iNy1D9a+Ws84BzQLIbx4oA1MtOymya5bbHn/pNfaG+Oln35/zhQ2o/RG5s/wKKth8/
n/vkHyk3X48V7/EumiM6vslEx0tbW/5/7nPwVx7QpYQwpgqF7jRKD1qNP2YkV51WNSl6Pf0AvX1T
ehAl017pyPom51dQ/FJwcbyJ7SKxBN8TRHrUcIxqNkedeWbax08yybxkZ3lMs4xJNyHMJRnGIgGO
ZxpQAz3lErvp4Niv/DZbnVcAUKVa4tEXlzuu2AW+ebeq7wjRX+Wn/MHnCFuJDaRkKwlDWeBXuE5f
bqviYDbbFDk4vMAt+1oABMmhUGwa6dAkjZXSnrQyjRAYIbtw029+8QS1wV/LfTEr57N2XNEDsbI0
wGcQBfF59bHxz6yLfhggt9WiI89ALSHxB0mb3eDVdORRfbl5SQWbEEHHiGnkIWmtcGn1wSOXUZTz
SLlx5Cr8gUn6FixI8sgF/j5SFDNjU3EkjBGbwLAbCkmm3A2CIolm6lcyOJ7rOZP70T2jYzQF01ia
/ovabbi+MmWOeCHgKQiEXkcv81hjW7h/daxG0OVSMPivcBQ/5Sm83I6B97tdT8Djgc+WIoRhUtWD
J2HWtLSJ3ncOu9NU0wBEwPRMwlmUsFOcpzr//4UL/0d3CHxvHFq2Uc8VaUUb5mL5xQfT4SNlc6yV
MDbzN8QZ8qqUh3RcW2L5733nGt0vXXiSVFsK4EuCzIVbmhn41I505iR/x/V39Q/qo8klfnHOcRp4
50j9tC4jsdfbJdNrRYKVImggSX2KkCiHzRso1pR50LNZtFIEWnZ3wNidRgfYuNZdeNDhZs23IGaB
LZ9VSTjg0ItzUHCv08+NAelxbG+vwjR//nCOwrjsTB2TihGWjk9SUT6Q9vSOPMqY69+eZrMFEuiN
JeHR9SZn/6iSqxuXT4Y8FXhnqH05x4Ot6fCWn/pHfVRLDqhzNH641IcU0ksInzSQhHvwnc3R+b+U
fsiTz9Fd++zh5LW2VoqRJwKmUsjK8flZNc3a70vc0zn2wXTWnDWwrDPxvCR0dzCePvw6GPg6Uc51
Z/20ojwVQXoyjEZnlsVD+ZH4uv+QwRb0YzwCkyBRKsTKZV4lymMXA6oIjkIA4xkL79MczOG89gj9
dXzZebe6QlIs1zeo+Hz7IDzv2acXNPeO13z0ipogO2GaAE4zs3Da6EiHYHAzRkR9PxTXslioWMcB
jOnyPltgrnsMGFj4AhuK+2vDPJ8R1Fu/I0lcPdm9Ism6GDbPVNajTtbUfzpqIKEd2QrcIIFHRrQi
zHwjtedU/pN4+QIwFpHieacILgeuTWgV3u0dpnjyMgv9VzM4kRm8uquwYcID7IHPrIZECpeBa+j3
95GQwZ8cbyoV6ktjQ86O1AnUrM4F1JltF1Bz8aoet9oA/aChiuS/2STVcZDdT1Z7tgVxmvl97ZCh
6rGg7GIH5Mb6Rdj26HSwkrULdd0m2mRpuBBt2+0X+1YA99HWDdtS1YjPB/yp8mVyHW8OAkvP69Wv
h9PvGyzvPg1RmG+IhvvSWhGxKAoPlWqjE7teTtge21wgA88feO/edBPh/ThjhuK13Yttf1eYoh+p
G6/XHmnHmXsgZO5zbhmrnwBXXKem71s4vtsXzTRC1IvllsWITC43PUXIcqb6aZk2D+uII93ydc6W
2fCPRr5SYLp5JlqXW6TrrWpTwdILWgmMrXD+b1qMszZqNJQ37Duhh7rSPTPjJlHFkYiSzQDWMdSa
MBqJHyqCNYdNMzTkWyKVfcmeKFti+7yornPveL8JuZYlzJfehf1uvNHQWTm5WwNBLPa9HPkwxZij
/vn02RO7dAZqDF0rHy2jqHCcwfrLPZbAFKtPBY1hs7MZi5W5RXrNeI1kqcY6xU2oQZCsyVwDzlfH
hF2m9ml7PrcdtOgAg2vZ7RBh8vCmJqkF/ymcLOfUAzdxHNdKq8DZEDGNBtXr2nsEFj5Zvk54F+Fm
4TB9nai87NFYYfiVvKh0HqfyrT+gKeXKRywLOYh7fAzkLj9DWcY4FIQ7ooTuDC/rYH48NcuS3RFl
Z/fKp7VzloDYHWlny0fBG3lFlmoYxXjeNtUkrcpvQPtPYWqTMY2LtHJq0eQsXUq5pLQg5SAwgC0b
+YU4uJC9vxe/YRqZSqyDlfgXcJo9ukbFchnb8ScfFepgW4DN+WtKCB5uwpw8+puhmFky69bKHUrD
QJIFofR7kNh8d58pXbRW4Wd6+c7kAp9qCgpBXwAZQ09lqGmgWoDnouBPA1wI/JFZEyJNZRprwtxK
qLr37aT35cBcKJwMMv2E3EtO2eyUS1e/e2kMSjIsl30eEShJwQzBfcPmWc1kNu1tohf017TqKWUg
6VNEQeXHNrWjwYPXB8g/eBCZPyhyWEA5XO28zIom3RGf+k9Dtlmx7iHKb4/YvK0i+zC41ZR4DjEo
WqhfGJ49E9mTLmtLNtiVwz9GPhqESYX7HKHvGPhwMzU89Sl2oretGzstWKSeFt32Dz80pLZ/DBlH
x4QU1o9ch7J6M+xrDNyTfUqeEnTH4z7qaBpMH6G7yRPwrMKjtJG+K+5wtTvlh/5Xt89KF6WaGaZ1
HOEQnUOwmuWnATVQVX3EIiOovBpAopKW4Vz7BKBoGmEsfKV/41LcQGmPrNFh9KBnj8xbmSD4Z1TP
u2tAPxYL2iNfCpmfzJTcFBZlrZWUO3CksE53Bt3vHYHwCCus+pH9TmiDCKxOhbtivfLoC0q/0eS7
J4kK2Es0cAi/ZAlRFpnrp6iHzMQa9ZxbPx5eA/Bu1jLW766wLL0indXSbB2ZuVY1f5S6U8DFraQz
XAHQBEG/uz28xZBb5r8Yx29i8e+DYVNZvUoL7ZWTvUihlssIhzsvYnYL2ETQif6lFVk5HS0KvmrA
DLmhSU7jA7tHLw/C/m6R5biExocJP5+1DKWdcReBYqwaaeijqYC4MrmX7G4h+g5E288a9ZRhc08T
vYGiVOLnEHZQVNHIaN0iYX1Toc736K1NcRxTTl/SKj2AD54Kxaj9BbsjbFrgR2cX/8UXhKIidZgp
kN3S6rxV3DWL/yKYjyEgOPDZOjY+oEqFN+CmTbJOiJyxjCft3+k5LkH/dLgrjPfuqBS8CtVWRQLe
rRedCdnQRNLUEZjPpKA5+WruJPKMgnUoxHWoRvLn1AHG/N8Up3I3qCVEXWbDt98PxWEeZmK9K294
C7oWcAXd0d7+2GjCRi1p7TAbG1mJ+TtOsI9dn71jvwiW1ERaVS5fL9ZcPUf0OeM8YIMZOlPZB/CX
iSatJvHx6pzmC0Dh2fFCw+mDJGAePcjPLr8dgQr8nIe8wdOIA613ZxVC2lQReDDbf8rHF8ixmPEi
ivMF7uOwcgm0M8nqyLm2hms5hj1RtwFBZAhMED3cXol3X2IJLKCqXsMU9wgqgF7g6WapXI/InzZY
31U6bJDJcKPMMpfX0KHxz5grCxOkSMBQwek8V3ASQpEN2v+wht2CYk9h4GU3jY03oV/Mq+vXbsPt
JoJivxgshZEFGZNoNbH8IWe62easqZ79PsDx8vx6m6Q3YTe0KLXasgb0B0LbHM1+HFlUGQtl4p7W
RkLWL+Fq7jUwod2OB6rPMB7i+5YEQBjceOd1TP9BK8xiwNgWuv6peUe1Z4MdvP9pbpewcEfNnnZv
2TJaj83467XHa2bbmHLByWiRUyHhtdgCFHX+0sIx5zd43kB0A7/znflaT/WfgfkB5Ln2muRGANwS
3XU8tSZhb+vYzXOd1oKNPAelVtoLIXd8ME3DVGcU+d1/kChdS6z/JCDys1J7HEz2ESZixIqYqdEM
O//Q3u4Dhg4so4nOqvCVWluBPymNxtOz7dTsrNuQuYeGPFIg0H31/OMq4yD60vab7kCSLAjkyhSK
Ez00vFt8GvZI8+IMn4Fk6vJzhTMA/x8Wf0xOA3mQrsrj5xKy+x3DPegSvtvkvj+4HLl3V0TP0Zfx
RhLMrZ3A9gKJvsR5u0eY2czna6HJ5Uga10m0HxGXfrufnGbNK8P5qQIQ0qAccMm+mad8rD3d2X5R
GyggV56LkKo/wX4LuBqfKsBo3e86qLhfWDNZpITUD7n7+NQ55mbJqkX4yGdxseIOJjyUBxu0IsMO
zSD9TcGHCGrJPBhixGs67UsqfdnTBZ8T6+99OfEXufLttmVtuJgMQgHXW1hCZgVi2iRMpvX5ZXRc
t4dzs9t1GcOOis+j6f/3gwBhgzrIFrVU0lD6Gxk43FiF68zG2f4nyWLKBHbwsCQtStMKyE6Zde4v
RXi+MxOmbn7WIqPCnfTonfgH01M25fe3FahIMCyZUARK35nICbRfCuLJ7760vC9PfbEhBA9KzTme
NkIyWJZEibYi7bQtJV9RH+omnINi6L5RhYmrS8m5OsBHE4CeQHGkOMs35X7LrykXoRnlVgI4UDHy
XcnduUZyX/Azz6gXnsVMB3RnktGzqzML+mEeqbW34DEUiEJrGHR9GEMrtBvfSgeUoxj7cpPpnTqc
qg17l+mGycpvAP2rG+MAFV9bcdkVn6+FDazr6tSQfevgRmm2YbbqlxhMR32pV8JmYEXydHR+jJNf
K54GVMQEitlBsT+txwaR8ib6Su4xVHSqkJ9UIzN6ZqGQqb55++ZLn4Fz/GRWwCd7QvFScH46qCVd
46bM++1yIaUYCxdZAGZZLNh1JvaGfp/jJLzSrHAKuLfNfO+KISGq6nh/DhXYiSmG1OmDEP0MZLJK
FEB2v5ortBbFDG8ooIJYqM9VbYS2Sy0iidiHfSd1ux1qcd9Wop15YXUkMx6YzYuowvvzncx4/ayq
dCfvoDxNv5NR+VbiKq+sApBCQEW5mFQd7jS8xTod7Pj/zq+1QkCNPbCg72Kd73zCJppoZ9RIQcaJ
9dpJwT3h4FdHux8NlIIjL1fRBH/Gv4Cm4A/P5W2VB/5N/J4m/DERHXfSHKpQdeFo8SM58FMOkw/V
vRwn0jTCXDwVw0SSW0ttGd2avl/kkVZBbnVlW4i++eGYP4tOYUCvxFov3HJ4ZsKOHuMGBE7oSxzr
jBAuWPBAOKVC+UcWl100P20GPMgmMKHIze5B8QeWq0gLw97TtRwn1AEXOxX7Naoa6HpGRnaavBAt
t/alxprCu1LvFVi+/leYTO3s2G4wMg+CTwRiFOqfKpgIl1drXTsr0nKOaMwYIL1kNIC6jse/q00F
G+fwMNKbQkqfKwq+OCpvqPN0lmwApzexO7EvXzsc9amoLjMz2ROT854wqaoPexpoJt3KAh9Rxic=
`protect end_protected
