`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R+TTV2BAhe9Ek8IveLCAIK+vyB2qa4TorazWyGCbrxCKkVhTBvAD6RqPeP/JqtRuh2zDPzraR9rT
gUyNSWD83A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XM2mYTm+gCT0AhW4S5p7IlzH34WHm/fa2tLSENK5xQp44huwLBqk+dBcYbe4GM+6wqA3pzoUNE9T
SluI3P6DpsOt14ispiaJSciB+VdlU+Q0e63sKyfq++TGO3CTW5OhLIxojUbYrTbdY4WbGkk4yG0Y
qGwauBBx1uBueCA2GC4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
M9U+BjMD5E96pT2zTDB1OSiHn8IS+G+aDNa3MIF/jeClLSPAOJwufjuzRcyAtwx0354Pb7AaFOwR
6CcoWPQM1dcUC6avyG/0PRrtZP/KpXS3/9PiWsaFHPYVLfqBMCUDoraXwfpfMxmOy8hD0iI6TtWc
j1xJUXVsbv+kqOeTUloYmwdRx/8cs46FvZfnFpiZXMFMsTsT9zvmCyNxiZefgFKT064BWsCkg2fa
W2IXperFJQzpE9mXVwGSjl6xDUp55esPyEPcDI4xy0T+q2KtBQj2Qn2DJRZ8DKAvjXNQmo/tbweh
l+RGgbFge035kxDZ/t5pFweR/SYowAMdG2yOwA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
absLoVdCG0/WeiZ9M4NtAUjz+XnLze4vahkoVw40DL65GHoB/ikdBh+LyLQ7V3LckxaJp7Ihe1ow
2yXZZfuygvynBc+n/CI1EDwjo64cUTgVLg6gqySahs3D5Xkp8kFBBxARQmdoErJqqhefej6SXrxx
13OxNfq4vRGx7YG4l2M61gUhVtUX9poQdq5dxitmrLXD1kpdnUsj/YIpVBaLv/TBn9G44WiyRNIK
ojx9q2JyYKiWBfcBh+fpJV9PudrBUPMu8kvWsRizFr+r8Ya09D3o9iJUZ6FWOBiFsidvZNgmp1u/
nv56cp+qpaTesLtwmKiZbrhQtq6YXQvzPpDQXQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
t2oJ825g01R4DfbjT3g+VDPmL9PAyVC2t8Ozl94Xb2xucD77bNiPcvutyZFkA0lqWfRMp8Z3kkTE
OOo/FpGS3c1SP04/jMKLZD9E7DL6iVBRfxa3itPHxsSD0RAP4yPHw3yCiIsmB0q25x8+so3h/QOv
DKZh98m5ku9UnG+pY6c=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
koDeaCPE+GNu9rMKu+nnX8UvNKbOa7mKCRwRUXCmZNo0yL7JuxnKQiStr89+6Ws9bOIbY8P6XKLC
WoSokcQl2MIZuh7gUJ+LQSPTB9HIkHPuGGPibAaiYY3e/6TBvv0+QG5gTvuf18Nz0UQyxRzNBFY7
2e0fNw+zoh4XJubbVaqqBBqTNyIM/naqx2G+DBhvJF/RlcpsJUe2eVt+uttis5ukRD1ndenp7rvA
+Ub6MDtoxunfFJsXEQ8QZkuZiT5XfcmJdkquGywSafJqKksYNJZpGleQnak/ePqKq8cYIbfpqOo1
MlqTFX2khe/WU/cqsW+5jXmRAgWueTOvg5hW2A==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wZaMVki09KtetQFaQKbOEpc8bkgxHSc8zyuzh+dwZ44uN2hbx3K7ITnC8dDkn3EMZGwk7C0u4eBt
eru14n5jQ1LfuUg4cKuwRNAgFxc7GaymqPYSRK9OQZHWZ+w6Alh4X9YWb6UVcsv4sCJA8YT9QeZ2
8PJYA3L+OY2t8Dcx3JcdLeVgMWDrP/zfpXyfMdPpwgBSSCqJHFsYdlG06onoQq2DDJ/SpC0W2oHU
JJAOTss7Cf3giWx2XTrorU5k4KbClTaEv4QAsogatkMf+oa9OfJQg5b7OUNbNqSzTV2IvRXtKIBC
N3mFkAtau93JXZzbow8bF+Y708RmUyIR5AX9og==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gidhQdKtgCKZpycO58SKONz/x64JxoYiDvm7CY7FhAgR8N3zqVR49qh/d9ImLGjAjXhz9ISSvhiE
1TpzIsqbVIoSEHhHCsw8fW3eNfjSKG9+5c0qMghoZBwnf9txWcso6wczPV8wSYfFgOnId+/H4w2u
MtSdrp2j2HeGCN7hmduXDeRIcLF+ekxNNZVk0wscD3yxYdFDWscebLgM1N+Cx8uwWvloVVe1fNSl
IBecuxue/tBnCdqw10D1fC8gGorhdNUhO2bTYqZL/+voIIAXkux7Z0BGx6B2uSJYuZ0j2LS23yyk
r0QDrL3YOpbEPBbFhTy9LQz59rkITBRhVeBqVg==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lv7TtlI9EkMH+4ifu40NSGcF5VLP+fQr0uBXzvHjgpvggoEPEBlbTyXFtewlIbLNuHO4GjqSxFa3
oGjcKGgjJ4JKEHh9NZ/42sDCCnN1TS1zrfhPhpg3aJ3aGsOq5GxB6oAuNGvsTC7HgKk9lvgZfAiC
9ubfhd8fCUCrbS2jYuGLkpNxtwRxEbxLfMa6l2yusSJt8g6sfH0aGGBJWZjKnUZ1SyA1DmzZW3ox
o1AE17uwesEX5+JGPaqlsN+jLpbHhpv24GF4NS806LjJrXOO9qXbZScc78Z/R2xMBhLYAC0AHR8o
o8hlz9kYq3NSGSCdEMOcxNjVxDMYBrdZ+Lc+ag==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296400)
`protect data_block
ZTZwWwc9Z842HL5KhwLwFSCMsopuB7FReqmWRPca0chWkSV+hfkN/mv3fj6VpOi9lLHydvcR0mAK
xFpmRBDXwQNKNOJO8WRztyVw+nYxvKIZspNGm101g4jQwG8TnbWV0PXzOfekM6MmPNRvIPmXNAnC
b8t35pbRwt82GAQHrwQhlMeIDbfpggpD8Otq1T031ptEtIu9cknB+m69RCT7OlRb0ns9cYJjENwI
xIVScU1v+rtsZ2sqNVLeRnykypg7FC37thkYVsq3o70tBLdtwfSq0hHcBupmEg3NHu4AvaiCkech
Fhz5+kcQHutHPWELvlo/QQnWTMwkDvnvm13BvMUlKEBLJVgZH2oRK+uv77ZJlcGdB3NefgSJE4YO
aCc7jDVqVYWzlDC1rXsF5CEUcOoZabovks7YRBc4MuSoPDWUbbQqQg8Z0/IwVP+GooPBCMaWGnM3
55oJyhPznr7bLbqS23Kbw/u2sV5YqXjN1CnybMrzozMLNsZXkzQqr3VVn80dyGoMe4dC9ebuxhkF
WHM69mfIlCG1hDgC7p3x9+30lutUjM0AbIkGy/P09/aBf7VuDz+cHhL62BGrGsSSIQk3L7yv467w
PRVmaYE0PhsHZoYEXKDYlRtTdjo0USw8FCdOhXis1ZwTiLI98eptYbq507fqAl4u79G6EaRCGce8
mx/10EhXHeFK+9ITDDusjM9A0LfOWJOVYLA3eirG1OiqZ6Myc6qeIY0yaw5jX7hbXsR0G4EEvxLh
8uHtO5yzuJfdFQu309PL8TpTI4Sywy5ItLCPLhbNzOI7V58DKWTjuSN7rHMEDOiHPJcDDkRwM0Wv
yOgTc41bhJHvcMPceQYPpTCwUH++kbLUU3ppaWpHhMZr/CNRCdZNWcM7oEgAX3G74UbfkBTUumcf
BeqzVPwPn7Sy4G1+TPt2Y1mzmLQaNhiG3ZOC6QLB5AAu5RAF+RcY7kX2XGOYucOUJehTdaY1RW/S
ecpBuvVWIBMe4gsJ++7fYlaDj+ExDDXVYMWt2bZ4qm1BndPxKAq/ey+MA8UKLxJJr0PQHj9+bZZG
+lnXkxSUw3pZUw9CerY4c0uyNGaKimYc9iPpzZRhmXaNs6M1gANuGsKFe2ui1jIvuHSKgpqHkrPQ
fN+O73gYZbOPhAWlkPJu6brCvq1UWy1DjmDvRzwk6WRBCd4dZrf+YL5jOkKtmJDGgsuTPt8m/lya
FLkBOFuL5D4mZLcqZUPdB0kEJ29SUnSncYmAxShJ5Zx8Xsc5hv2o+71DhPaS8gN7CchGqU8yLey1
O9251qfxMIWGe4r2KPeRoAg9ZwG5evNXZdHuIuMS8zTHlt/vniG0NwliDIaGW2kDoSy4/c23w2Az
v4YF8VhIpUQ7iqdf3ZdiD5yASIm9IwL4QL4TG7KghuMwD5ZMavR/Ib6oSbK/69CwLK14BOohFXeB
qhFBc86RP6xqFV5zl9QKrm54rOZ6rIlRFjMnmOxZuCzC065ppwMiZijL5vQ0UCnH/h/Q/Kdhpqxe
pQZ8XkdMmWk4CviOGErVXe/5SOgMGCqytuh52NgO1QUKj4PriKRHvgUWwhYMzWri5M18iEJ1pfdu
JTHbemkxPZ7SMMaenH/oz7To9jioyZbJIYYvv17MSs7T02Dro11prTPB+ndnkIr01xiwym77YHAR
Ek7rt56+VOBtNL77yyWqnpyaBN9VjkWGQSWCOGxA0rSu3m/fh3qSzLUGVqL5VuRWBrZpvRPahjkl
1jqAe1pUbS/NUV7JaUWeHqJ06e08L/f0UHIrb9Ca3WB4xTUxPTEtsofT2SUNUHJ7K1gtYk+3nlQ0
oKOznXKD3LyNL+74s0bXAhtzvX4R7WbvXyVIKhly1rDN/Prw5WqbJ4p06JVn8KPn0pTZn+MUSRfX
irdHhfed/J7e4N8HaRnl33P06AnJ4++ypDaYWTuxvXqiQJhhIrL3i4u6sp69QVLBvvVAG4ymlhp4
p0wJFSur+ecqHTqDxjJCPMk0g//cwTYi1iItxLLLIFcMcmqIJPwlssOsWekHP3pgJciqfpiqVMsJ
VZNxGhn7KFhF3c+dJwcpP+EIMOZ5Zr5JcbYaJ1mOtTvBOEcUXE/bsAEo8VTwgQ+Pq1Q/GOCF12eY
A8q0E5zpamzB3fv59PORuUICvXhgrnPuqCgvuvpIJ4GFbo9AK9zn1TE8pROEev8dGqzU5JbMdcli
Ku9Kv6oZif/vYjJ6ieeTaVyThNuJpmyit5iqCW4sCXAQJU2IicRNEi7Ixd1IpMrvkw4Ciq1GmXfv
wP1u0L1WfRqGg/VA2Lmg56ZUxHzIYgpKhY9UurHCxOM40sl6/u8nCtuGCu5Tf3T18SLRVj+obMHu
t/9REppnoNb/YQwJ3hpeKLe55HEWr+RkwEsmwJX67rrpghv81NQJkxo+VLTjh3K+Q4Xe+bEmeORq
jPRR6vKJBqy0w78WDRqT+dg57VcGvFhVq2b1dSXY5/xsVk6Ntpq/DALB7npC4udr2eJ7THKZrBdR
VYQ1jnSPXuunZ171UxEex2ZwStqixeAhx2OT6vz0+Wv+roi/GKlCM7yhRKr3sOiu0Fr0iF07PzDq
nhiO4K09KrMpuHoUPX8TICXQqCvdxYkUI2Sh2dkHy6uV/DKgsYewpkENCbFsITJqHKfLlA3Vpg71
zzwyja7Vy4FrHI0IHTFS/msoQkAuhPN556E/5kf/Com/1OzoiAQQvoVmXoWW4TUxmDf/+dlSasSI
QC1qC/CCtBgUYRxmXtSXRwFHVRQQWgxyrRrGSd9IpgS9hviVM3Fl901rWzgaw47R7JiSk5RVkWYN
IWnp17EKsI4I5J9vgScuI3XcNo/Ql3qFQn3RMLfOWlVHXKvQjFHhtlkR5XnxG+Uf/dlbedzJb0zR
ExwyQFh/lmrs9a5D2VZf8pY9c2eEFtICKKW/jMgNvxFxw0+uJn9puj7qeRtaZ/tE9GYQ69GaimDt
S0w0RZFFtir8kvJa/pNODXMYt6fsWXUPuVQLhk+lUE1abyrbfQcuWGxbVzEIdRx2hqACkwelknFZ
jbQdBzUngji9xaUe/Xd+yKc8X0UPeItXW+fclBk65KwRhU7+xllSJqEfmr7kkQg5Ee6PQNm6N9W1
pDI1a9x8qa6hy3xBx1OW39E34wuT1GVKKb+n46TCTf4Kbt3UOW/Jg1lJFey/xOqy2GD6opriEYJ5
4t+NXX5MGZjDCH97QemVjjQB2Luxq8Y8px8m4RmN0tBGk4I3+hZMEQ8TwjMyj2usGQgz1kmdQXSA
UINH+YtEAlohjl+hBQxCv7wAIb14MewgZDoMtLPLZhUO7yOSZhHniBSKbh46Ew5cGl7EbGFFXicp
hy4nwNlUyF5OBs6YKKx83n9g5rUAcgmxfwbeUeVxAoNRtankihR9zNp1NTyoDXFD3bGXTnXl3ueE
ewaGbgPCs+YTIaecZNlqVKkhdjDMyQ0MHSBku2z7a+H/O1b6JFyGKhePmssSTWbW2xosOW2m9xo3
5arqwkg6bQnwLhY/k/dSQ7avG+Cax7n/gXCNXlUKGfYIsrEbJhFVeVibrB8eyLOiQmMu2aB+NyZ5
JwKy59wS+Z4LNZCQ/tpft0XTz2H3cf670kAeOaaHh/jMo/gaFwj6IcnKUyeDojosbrYLSq4ekXaU
Rxe2hq+bdmCiz5c5W74qtjwrEmYSQBmfbLiNwTbN2LBd9XjInvifsAuN3F0h64mQcUyyamFMBvFj
ijAiYnluV9yxSQ2HRKXlzfqos2WypLK4ZufbpXQBOePqvrtubf613GHFuBMl36BFrN9Z0kZnRK4M
CV//XN8KlTzMMDE1Tsgckks96+OHj+f0cZwoyMYx/J0OMQDa1UNp5vWB31qfMmT5Dt4pFhd9wlCH
fk1+52UcFPfwRzq/GvvANW3D+Lh2lMV0N2M0BAtY6ioSZ6EcZUewln3e8vNEqd2NbeSsAlUxHQR7
pZaSn69+BugbvRsY2gxJWIxfp/AdaNGJI89jzurCXAgxoOdHhJLmyo71M8gC4ptJo3v3gKzV960k
jmaqYMnoogoPssoNkjmxATbH8OsMT3P1VuAYCpWD/xV+3tR3oz+hbCilGGevPTBkAuDGICs9JcoU
avqOPuDT9VYaII4b9WjIIO9I3Upv7PxxSLDrAqFwkIVNsG8wDtlmO+0Av30lV3QzgYMbp1N9adHw
jDXPcrzFmm+x9Ct5rlwOnzpoT7ZOLC3brA20eRj0zRbfOAPMRJOtZ/gea8rebJ/3DB2z5Hrmvt4R
V6tsVJMqTPwGou54p8w9TPw3MbalXU1kg9ZQPymZHdNSpHv9Ur9lfaZRX2zId8p+qgAADsSAcwQG
5GHtscBM1T+CRioia1XtyXe8x15crGkB2x08kR2OLYlDDEnwfG+DZnLoMXC6AulEk1UYJoxEMGm8
6+pmZtUAuehSBshnSO+0Ih0KNpara81rVznE/La3Ywz+fROAvE4D0MYHQ3oaaWav023Zhe2UDKo5
+hBNgtP4+tkF/llQ3ji0yNhYYrI1AH7rMq5cKHJOl5BD7LWSLgbhL3Kmj1tEKwkAXGDij2vf92QU
LPANHRKgqpNuYE9y6U5YGkSvQFRtV6Is9aMLZKh/ScsC8DSQd8nMCUrZ4tcEYAhopQfnOWYvkYbS
gMN23AiyqStol2C4RDI77LbIkkFYBtVM40Knh6aijEsQBQhyS1ARksuLcbLwZ35/2RlwMbjHwacE
1uZbKTQjGnA1VkHZy1clZpH3TIlyLUgvxaGEvNLJLZ9N3/D+jXjWcjTqjjE3yxUVHp+mBZnPVCpA
4MLG17+voxI7fQNcKrJhRqaCFMCSxxGtn9xwbWNEWuVcGmVaJOFg9iz0d4RA4+6b1eRUIcw1NP16
oiv2rkc59vfhsvK5kAm+3kfWstpwk7npwl30FDsLWFIg8NLhfqI9sSt0qfphmPDmotQQmLKsPTJi
uWQZsYw9OYrAzFesk97ibTPmDhrx04yBwgC8/U0qDKQHjoByXgumdIgkTb20rWyg+udDxWOX0oIA
IZeXrd08iY0XTYfimtPFPSFve8x/BXNbLIpXG4TTpCx82ean7Xx4IfjQ7YmapPOmwfDNTbN2XarY
QdO2za+PSeHsa1vS3xRyJvUVUV8ELVvFILuch8Gpx2vhgRnP5psS5e/690fRw7VRTUsIHcu3qKwO
V76FnlwfQpwt7ORS5VVbrkwURb6wvLBP+n/Sj2pMGZD2ymizNviJGA6yEz3m0hOCCAGKVRCCLzm1
CkNoHRlnuIzwm7LC4V9SQeDg0tXn0v10yVG2xKNmBGoiaYV8s3Sivo0aTWJnKLZFjj2wD66CrpOJ
amuJlcdiwT2Q4E6ally2WGeSyy+nPG9I8ZaxOND2KyegDGyyTgxIeCqf+PUbMmR3YtO76Aqbv4oC
E4/nlu3WSF5rL3Y+upRiS2qz+//Hh96hN5LqZYVJ13NMGRedTwivp2kdt/YN2EtIfThUOAfZ3DZZ
g/TRtxJ7bAl95CxD1k8u5eLbx4orom4cli/WRzq6bjuWd7qQn8eOnMbwprHaHwAjiUohz9pwbQyB
9rWoacx9DSvjOV169Vx/dKaVZubhaRK6jwGvQ5uo5wQ9EtbiWIO8XCcVyDug80EFP4i9a+2wdOuB
N5k+SR6UeM1AvSBIEFHnbiiIKaoBvj8L4ZEVsh0Cw7KglhdU45lAxm9Du7mZWuju1GZ3VV0pGmEK
mG2RW7a3LRtKRKWrfvQdVQR6v6gHQmYF7juG1hkPgameP4GOgUKT/tQWkRSO9Jej0zzX32MeYOKN
6/+hK09nO1pW7d10jRxQZPSdUc0SLfDtIDuZ8WHHps3y4iLaMauSUNY4+8MAoQnWj4NFML1M4Isg
7SU4KpIZWb4MvrmW+8/1FL4ZZw6gdO1/aY53UxJJRxufK0i1zWRYd25MOt10rv6jJmMeypYx8ptG
GrQzIPqgjjrvRgjLPAupbWgloYKD7itKAsS7Tr+fdp/kgCG9Mk26/fJj+e1rWvlmdIeo/6bXsG/v
pzH5F/vMNvWWQJ881bDwQHit+bQVLT9q8sWkVOl1O6BZpnmDqLOef70vpW4UH3STMbwzO0NUA61S
RZ7jJls91tg+ar7CixzEldsWNSOcghbJCJckdK78iNsDdKGUxiXCj+Z5Z9Fj8q/iHNErxScgvGqO
oDvr4rzAsmbOI5q0DyOL8FLo/uWwK3i3K+SYXywiSIrjNeZztTZTxlAcyNk3YlmcDwpvtgYvdwdg
iKsIlnXTHPIZ0FWfKHDkcZN2i5hRuGAkxpBjbyOyoTRY6jf+KeOkQdh6HmqdidsYcl/fHzbXSzse
uxQIMH789avQlNtQrKC87CcvV5AtOhILGUWME+/Tps9aVaci3qvjXDSkR+y0G2/sWJQgWiwnAlsv
Syx1zUwT+2Z8xuxiQmwvzIbkNlE64GE93tMMPCL93626rcZRYcik2YY4irMpETxRVWg/3Rk5cQCv
f+XpZnCSBd5YV8qbz1dPo1blizSp4elJEwch8dxlzBc6WjfC/VzTK46Lujy+QV7YBrr8giwmB90x
S0oUAbxVQrUb72awIq9YDxsO63eU15CpX+p0xnntkf4Fg5sjFLaz2roPKMGL15X+2GZxtVuuqjRA
bjKAl8QrXVm/U553cGHxSNsuf5O3WIlJiFXn/3BdPeyvGqOxFqIlFAWu1/bxKXPjG33G41kvSw84
w+WelQ3wB3nizajRn0wkp5YzXTiLpiNosm7/9s8gzRD95tTjTcLga35DBjrcvhFNZt2KdO6StcK/
qFbF6mWXnLrDK3k2PcAkImf4A4iwvCppLdJxTgE88yEphJ9scv0PpjUhh1TfkFJTn4f054M+zqvT
RaWHafzjHNNSz/LcrXyHJaYuvDc8uqE8aZUuNa9dQEVaeudj/6Gk/qBzjRSWUWnZboJh1dMmMtJT
nqc/tOie7xWW/nKT6cQkxcDcAHVeFEd26wtOm3PmA2n48zcCvGKpsPNvIT9rvbQRh6X8n0+cOMcP
Lol6boM7LUUWKmH7UsR5pLFssX1yZ7A1yCYIwUoTSdCRxgjRgT7L0lh/jjU8T8XS4dnjR3QhTx7O
ljoo4mwHA2iejve9dxHibIg3hkzwwVxgsOMLnrA8OT2JounrcSq9cAbKZ6lFIY2BfNe8pe0eljqj
tUkCi6vIJCyQa8ujxwXbPxRskl7s2mWNcurreXY+lfBaUCQ9B0bzQGe7aoMLfuxOdiAXyIM7tacQ
eRA5Hxcw7CREZoq1LxSOTwYen2xlWcyCZCYYy/oTDP03Ufua6R1YSqIIkcxL7KOvB+rVZ6/zJdle
q+21YkUelVxDQua7WYm0TEBkEo2AyNuhjJP/BFRq5TKeBSzw/JNO2DtWi5Xf6fAujuw6VWsUAePu
vx/6DV97dukx/Krq89DRGzx3t0zd7s6ha8fYH4gUQhjOXWkMXr1/Ymdl8nl1F95r7JgyuksfHCom
eEnMamhkyuEm2jM0ateQc1KpN4YoN3HBHG6CKjZT1z4Vc+wPGmZoITarBak/16cTT8K1eZKKRo/t
mZZ4WuxRJAjPtE83Ze2qahLmuedbTLSNIesG6/fhRpYpUE9WnBLjXscTxu1t0Vg77AzR0LXQ6+KJ
t46ZZtV8HH/pHIwtS1k1C9RQNZsHK+Y+UQgoPikPpA/uL7r0QwEZv8U6sNUcSOm3VfEDP6gN+L8g
LFUoZ8pDlcSn/W10njuatB5cS6AERzu6pSCyHRThXOF4wXqtnAFD1j+e+ilh9W4PZKXHzIl4vzsr
8OPHGzwokVdfQgcMpwk6koOux92ewACOqKyXv9T0T4LaeIH0groY++t3BWXo+tF8W7/U6MQ8kRZU
OKwbLvuqgvYWxixQq7nO1OfxPz3QqdNYujsx95P5jDcweQ7kIp8EhVIq3KK9D65Ay1CBRI75teRc
H4z+xLW56yJjKBaPI3DsnxeRozWFMFCCLEFp4zrHnGHNpkaPkwb/U7/WBVaQsMqrfss8NAk+mmo1
pExoj6Zo9iPhPgMrDgZUubYMFVa3WyfY4897RqmeYBTp5ICPuwdqoyvcbXG7tDwxxoXDSEonoIgz
A13B29nw5OnhMHpNa9jc9dLiKmZKeqA8cYPIDPhG/6SVm1YaB/AundgeeueULnlyrPSd6ia+tyan
3DLlsoMzYFavP69Ajwo5mCloihSL13l1PpxDqLZU/M8Vs7eLMT0Sybg9HfUU6Fquri7YhDB3XnVu
7CLrjHe6QpWClnLVC44mNGjWXAo5We/Xb8oUa07NalBFDGoJMVfGzA/LX/5x4Ox5tkTj+TOS8kiO
sPFHvna2i2Q5s8ik3IUdLmwdZXN9NOvVgId3LsTUk8iv0cqL8gI3qhbs8NhM90qlCLDhXvKY/llw
WgJMujPlZDnvaPBzRYJaL2xEVk9aCE5zuJFbPrtM22Y9Djgcug/BAwO8So15KRhEc5QdOyQWtlQc
GAVzwB2PAf712wX/KORf6U2j0MGfcpowx9RMBuc5W9hbAxQd/82vLiPs5ZzumW+b9xI03BU48S33
oN3Tvq/5WNJA9WQ7OchM02EyyTLtoaZDvlBPdQLqtBgS+Ks58e2GXF4ULvJzMhetuGhtlp5CamGs
mnjuNUZ8uZKYi1PyuwtAgPCx7sKuIMPK50zPIPwU9xKv1GryKli2VZ3y8YP5Yf8TRysdKsVr3l/m
22cFF0IIbGnVc2voiiH8EhzdfwfebJ66rM2g1V//rCiqt5g48BJkrGJod7EIqx99wWfOlI6bPAl1
iD6wuEuAbRSDOdZIc0+WIC8ZnTzvMtMY9Nu/Z/ySmFR19Hvl/OIR2mfF3W/dOSBO5yem/33YrXrZ
CcaLulRqBGm2XLZtcxeg/9uI++EyZu1znbviCESje1iH1nocp9Fh5GkpAcWmnwugb7Q8k3YFa/tU
kJ0rMlK4FHE4pN5H2DjKjgrN34M2Inr7PRvGF7ObOm6gNPmlORpW131t36U+L7C7t5Afkrr6GcGc
fJh6qqz8JEq9Cc0x3s0kwS7wqbrsmMSEdG79ZBEeNDMOyDoHvGKuCiGCaruHZ8iTVrZrgdCAhg5i
EyWWAGVZkOniDnMbAuMZuZFDVPVbdt/aeW03dwAS/PaHEYZt/nBXaRay5TIRUDMxzZ0krqZpzT9/
BctuhqMSGcIf0utCCxjQD8t5Y6uw7trZrcLI+RWmrX3EDoL2o5mhPbLp5/qGlLa0yYwWMRIHGx+x
aI6mLA+WAtuRjcm/3a+Is9JC2MsnKYkT6lGoSWs8lCXnvvouymbzlTnzwt+3nVC7CUsHfUmQdTwk
VUB4QPr3r+E1sz86OIcME5Tr1QgBs507HaEZjDWrCDJf481uVHKfFVD0AxkeyMlYWwY6yNBK6+Ea
oFe/2RaHLv9Rk2A69Or5ZSqSYnSUEMsn4FTKOsskNzXkBWPXgODBB5veFXXtpJ126zubOpuHnnG0
7rptQmVgr0Pm9lg/BSicBaeEGZtQQJOCb4Xq/cTboUtQsDrZW01o0eofRzDEKlwKEI3959nx4KEd
lC80ewAt0uIn/juAhqvxum6+oFAACDQcpepdTna1yx5HZZ4nq/ejRGJs9bAFHzFeohK8nmCHTl5q
7xo1/o0jortqjB5bSNLdZBlyxpf4Zvj9txS3KfDxz5GEfnbZNmjfAjE/0O0T9rg6K3GXgimie9HV
iTueFiukxAAR6BMzbgW6RB8ZVDjsp/j18Rtn/yFCr5UfrezqgRrWBjVvUl29g6P+cx0PIpjp1AB4
GO9tklaisuWU2NaB3TcLw4zapLy6U85jcloEGVSfwygmdntQ3Fv2cTyLt2rm0wjGDBSLEv+guhOl
EkzfLt9TxcPjcBVVtqDwmjtDKc/AyqV06r5rssA/b2LpKvozI5Gn5MIk7GcjQR2GGZpsq9BjRcuP
aILN3dqMNs1oyoeRFHrfrD+A4C/F5295pfQ0a+hv8CkmSqhN2XnL8w1snKaGn8ql54wWbeAY7wWF
T+RptgY5W7Ekwqq4CjEgEXYvkuniqtmsZ5St8+upVcvYrDJI2B9ORF1v97DA0WlmQUkQ1scFXgMA
eAxdaoDq7iiXHyKdDW/Qgt2sbFWhLDxl3/LTp+Xn8R8bGgn4x3xVlJyjINyRqdN3Wl5qYnOtONfu
Fmtv984atN8bB7QT6IhIlQgpXQsHlVPaHPYh+3+FshqfBXrlUJ6PNLLq41DSC2gypyv/ewQWW989
y+OkyERjyERaZs6TsRddZyhxMqm161kKl1+x7IqISJ4TUX2dPPXMwBhG/QoBAxBNuMEpWRx2JGuk
kqoabS6r/ND6lOTjcCGUmmilyFF76263UCADKX6MAluPPvhJIkRQhZf3y5q770DE/xFe1CKFiSCD
82if5MpU9iU9ByWXalDL79IQVyjKDdHAEjnZdMsjZWgkFbX5/Z9LuvnAmrP++QJvoKAKmutT9Yeh
YW5AWBv6Do75jqN93jwpxBVmbSnOATN9ckkWGSHi/1PkDgUwpKgxML1GojV8bUUSlmrwBhf+6PKL
coKwJlM3JvrBSkgoCrhChFmwDBlw8PS/uUMPa8bc5qLH3Aik1P8tvr5g6AfgsI6oZxLKPV1Ppap6
wG+JU/VgicDyVPg6sED/RtKOXF7Og8MKbV5Wh5Cq7MDSkNJUXktfdUvhaXa6armn71SzyeypP8Rw
3+1FSU6nlIIZpwIbP+zR96zBGAUPlc85HtPm31QoNSQC9jpiEzcEqlY+9AzFsy0Sf9x+PetBfpb6
AUtU6Hrf6C2ojjjeoS84U+pszxAPc8iL1R6oUC7GLnNHCxcyx9wds5qFKWD/QaOJ431ZWPO39BXQ
jLDQRrQmEDOtrUwGVtwsOqHYchjA5mMG+6KkJV0K+r4Yi8ZtD4DXmFbG30XqL8UkJF4+nYthcAQi
g1VBR6qgHCTkhKsAXrhWUNC+R/6yptD+2Uqw62FBQHCBQXXvZsQVSQ0Rv+jVrCsrkpJge7xUaP1v
uq95WKUTxSNyxhhkkUwVO/b9rgFaeobuB0/4HxT+jJSaHiALR888PS9doyIkalLLuT0kwUC5/QKR
MC903krRv3uyhV/X9xULCZlrTA9FtiqlB7iuAaS8MTWVd9yFTMzR5qXvjAbyKjU9mYlaCMstAYQW
GT+YuasBNR44ZSVZBYf8T/KeFyA5hqc/sWVP+oYgbHisceXUSxo1esj8LyMfv5MhEZ1Mll/iTpJS
6xvxONnlMh3TG/Fm6OrneKC1V0s5SIZHIlBlK1ZsGSJ5hEZohvxK5AgcubkbLUNPZ4aCXEHGbod+
62l/v/cxiCACIKaoHlz1+kaygL7XsEBkKIA3T4pWuD6vt5ODe6Ozn3jNCUqedkJZq/THj7H1D5DK
CPshccFxSlotilTi05YJBCdpoMq03YDWvKVKQtMv36ZINnoR7rp0o6bddxIX74UDTSPw2m2s9Qo8
U/a2IT6NajGQQRC1CHaVAbn5n18bp32BwM0WvP9Pj9Wi0gqbtk/EPVcCMjkTvG7Z4OGHzkFhVNrs
G+QCu/ZkoOqVJZW/8pzJ94eKxO1FUOAqK8ClFo2BCU4REJJovIIyNqriKY0B3uj6e290fwiSAHoc
45JqOX++VFqLplbXQsh3sBgEdDZ8TUV4SvK9L8iiRSujwq4TE55aizra0YggfQg13MvyTD/7xeAB
Z+kuR8E3A16GoHA+ReQSxjLN0LJx74ectRzzhrxdSTJMhY2bf5YQTy0yn/LDNtxfdTA12G88c2lf
BuQ/vlMnS3kyk0Ya0zwyx2X7TsavFJt0KejH+xCu6bAznJY5AGR0VdT/pEbohDnFUotcN4+wlQID
0bNiSg7/gWfxEjznNmEffRI1qbEYNRrlkvj+D/WLozly0MUEaGuBo7crsTKNdCkiVgY9HSxxo5Pb
EbRzNCobLMnSje42ZLicMYtlJzYlIwCq+m38tnm0fYFY7qQJrwCCAe4BAZpLjvyzsEzzrBC1Hzgp
2iUQnvOPqQUrZjBjt1I0R5/vq83Nd0p+UbYWp1fI8ftw70TvzcNwY3RB8zqEpjOMMOIPRDjfI0vS
wJA2nRFbOgajYEIZllurvt878fA9/2Dpe/YhfDxHwAJXRhdn8N9xTvRpAhak0SVvueWY+p45HI+k
l1K1+hdUcEXEofx0/myQW1H75X0/tNqaHgKVeIeS1Pwpa/n+HptXMwoN7XURuU0yZnIaNzyMwlcK
LcxRKOftmFV5OMUrLValRensfoxinCLuF0raf9ep86+m3XmuUIu8YvAAHocAlNaVSF0aPmGxksRC
fTfgQ7q/Gn0tSraipqWud7UdaczITRqueigVXKyEotwrRYvZYQ5YWbclCFYeUZ7/uKLPk2hE84mP
n1yM4GNcjbfPNyuSkC9rTcEWJ6frOc0AWYMe5v9voHFczpnND+aGYKP9L0gDoWdYAYJX9LIz2XLg
o/VlAXetVd7Zu189cbKfGWdmlXIiaq4FP4a3rk+msd93mDdTWBq4KfZ7jQwdgJuY0JmgETPVLgse
ElhicXysmCZscRbgyV5OJyo5koQ0jGcA7dAaYBF4GiSVYlwsb+nADV0VPrsYo252+PRhhTXC7J2T
2IS7iVeJvE+dk9cmBE9GohKVEURnAARjBd8uluF0LmVdJTdvhvYaGMzbiHUW8P2YqLu68Bo6B9t6
XIiTCuS3ZIOipDCRzZ1i6jfUo81aQ4/f8Zw+ajdG9hOJjFbKPtbkwWJM5XZhv4tWNUL+Dv8Ag5dV
8FP7UdgjJw0CqLS+vPr6O7iuSzhWJh+Horcglfz/zo5k1PEOGyttyB1lrBRihEjYUlNV4SETq1xt
vtu+7pJo27MOU57VlZ9hyD2Ehwj7sDkgNNWbKBVcjOhcJO3HwsLQC/oz8vypk43f/2T3Pdu7Y9Gg
F9S4VgwjmWF54LZZ1BS6wkat360JZKhjW+57iJKDOsofJXXhSBjny8oXrTYVmi1L+KUY7q3Hc2ET
p9zwl1dNEYcwcSrdbZDhl8RpTWGEinqSfbemq4WDwUti5b0qtDfKnrhkjGoJR11+HOVfm/7/t1y/
F0DfPUPWSAkuI8syyhx+22A5b4k7fJBrA72qGN+KC/P+ylVw7h5twlyP4K59MBLZaq3G2upAWS5q
X2lGwBuHLr0B+IzZMlIPIBtMS3d5hfMOT/4EZLNTcM7lW/DLSiaULo1BTG1n2Osgpq9R2gVju4PF
KXdCoRfbOwbDTvu0AUZTntryvwZmhx5qyUf7/YheOJFbWbsOxVWVsJI2xhE+AWx7fwHtqI9IE+uT
F+uouGdFNJ3/UHgRe4msZC7TPHZXOl1/RCNAfSOo5UaEfDjaUKM4X14Hzd13s9h2mDsWsk7+7r9i
e5S8O/6SbAzOX0mcPWlv0Wbb0egikZYl+R30Yb1Br3w6yox/Ip9TXoMLvnf+uoD7xgpufYlsti1E
6O5Ye7TJsejEwWOwVS73GGpQBk9sXtIgom74pz/zCQJKUxLQv2XPF9+0Tg2NPzcWdesyb4aeRefO
RPcBWZ/FOkvSmMb2I64f4bbbQnHoQvLWgiQnWxckjOwmDJENCPQK00ZTeAanmXG8miM2bN+9w6nn
nNjQiakcg1bRCS9qO2LE8FKlbk2zaAAlNBIkniiTSDRl/rtSA5W71AfxTgzRy2dqztCdKjKbEt0r
n9FkRw0jIHw//6X1PzFT6NAEXKdSq8FcNJPxHfhgfZSrYpVZwPshVSHHHQuiQ42zs1QTtc2D0l8G
wmP6Kem4uFwwGmk79+mHYnMG+if6NV4GOyV+rWQAD9vKxRECRnsjMYT005jpRn5ICR4vf/izitz2
jvuVupYXRNUiKxdIglp2ufAXIjNXRvp6aMlX634QGQ++MmpWOcih3dRg2DmSJvoIZrIiQZirRRHn
3YQs6VzhwmFcw8m/3yx9zkPKrv7HZXh49z7e0eWCsBTd+fcxZG9VC+/bETb3f2o9adzTIb/hTFk9
Xm6OrsxIkWvLYPbRHwcNpXFHkopSoyM4I/NnXGo+NOSNwCDJlfxaGIsTivFdusFt6xp6rLM8Iy+j
1eT7mh6PVJLU8jK9kn+ZnY330w55ue//y4ELC6X3sROFLXcMrHmLx40SduLDgN6nmRIjmIMVDQuk
l98q4x5MTUFLnfyVyf44ueV06N+BjDiYFMm7hYAvlGWhHgjNbi3Ze/bA0XaVzrhr7incNLkexA/C
1VTTkKwsUzO5fQG/62nWlV9WSzrX7+LGkWU/p5Zl9g4JFRmZbJOcGq6+2fE7ZiWTnV/BNBkFRN2h
AnhyMKkfFKc2Nct1DKN/84MMZzxI76oGf8z9RruSzX1ZetRWQ3yqYDqZRXqJ+lD1vhqOJcwr+hVL
TqdgzpEvgzsbq0h4+7uQIGCbkRmz0mXFzrLzBwtSRpg4CIKWITEEqiC3gsVfLrJXAvEfnx2tOCPf
pRZNXw0T4en5NoLiOo4ocUwOk+e5tXc32/H275JIvQz+5wBdgez5yUMFL3YRS0cz/K3LuFa4IFzA
KsBkqhdWaaRPW2Obyf//rvuc8as4xxipGk6UyZutda/Edigi0QQY2GdxVwECiPSYWcSGPFBUiLk5
tYNk9bKocSV5u2iItsJmzyvvETFvj2gYix68flaTz7GY0jo8NxgCl0wvrGXNEM4Zsy5bQiam+jb/
SWqVnJOEo6MfS46Zs8vSDJ10Wfm91ligm2Itl/AnIRHdPF55t+q2bUIsuwKxVT4hKAxgeoHVRBpC
CzUXj6Z/NnWvu11bSmT4BdNrb9E9xpbaB98m0q5bf4PCOuzktKnK9v3T16QywWzDOSf+AeudAOTy
8ZcgnM82/PBdITb6eLr5k9gotBG7culeOqyxKkvHm0hOkR2/JgS+EbqHmvAu1g1TyrW8+3DzALlP
pKVDn6fQYAvMBsQ8w6cU/ejNpuS3U1ztYzmR9msCnLYiHR9a3V/CnKwhZoMuscQpHXkZvrbpo687
pVdaSjuJdBjxgB/VhFAK4/TFI6MwKlZ8CAOw+ipG8yAfjSp18dVaa2omyhGUydToTD4d63XiF2MM
TBxBbVlf0p4GTzTiTzwU3YDeFaE/kUrRc3abS+b2aUvLR2oxCD6X5Fxh15JeQFmhGskcm0IqYnYz
ejwbJjg+fO6NoxopnvqgMiK0g9hJpfyw3Dod687+R3x5upK5K5qd2FSyAawYkRkj9wnNgSJ/ebH8
mHqt9dZ6nSCMtmcXoyLfuaUUYmqO8gBt59eYM7+m+tQh3nzcjGlv882RybIXydQBfRC4hiW8XPWX
qjjltd0Is+RsjdtuPngtGHRnCwzBBQ9LTPJChXUo+lRt66viZEEiE2AdbtoGocy7S8MqwV7+ShRn
7XJqehp4mrtDZCo1ub5M3Ge3F/MyZxxU/jkyA6uenlhKkwJ5kS9u0q7Y++Z2kLi0wXl2xQoV3bbm
Vg5lINGYedkfCYXiZCk5N1r1xWaMKEGq77U4LJD6cZ5O56XW0Vq3adK8ONqxQ8fOqOa3SjW1ZoTD
ahcSG8czgKEzF7WyspTwceO8L5Ox2VPOH6j+nIkYFVfNZP02dtwi+vwo4z6CQtvyrXaM/+XHaDZf
iFvKawDjYZf3S+v7SQOmVsam2MfTGYrr3Fo1Xs3bcuwE7/cxjmrrB3KhV1TYA6yN9uR/v7u4Yjiw
MOJjLfCaYSv/s+cDGoHRdCmUmPRQ39nTp5CwNSd+TNH6eIICW/tU8RAVvHyg0zHxlV52zoFzbwsQ
lOOBwUOm15AT1NrlZAfMx8UiIFlaJPCfcll+WrzYmTvdw+fcDydHa2TnkFRtnWxLR8UMrXig1tjx
QAqlj0oTzLLQidJ27NILdfGHKkCXOD7t8fDjA+SGpdzEIo8ZDplHgZHqUe4EUyir0/jVIZiypytn
GlFzAasFT+5kSmkVZy4HjiC8lwkzbdUUULbgSHxzi8d1wDlIBhavI2AjgqZqTs1fHfs4TPSVWbXE
dlS46WFxl4Pyo9t/KVMseJANNycDWM2z6amAoXp2TpI8aNMbSawLU6ih8p/uUxz1bF1bh2azLCSf
+6o75NZpMkCvEyX24tv9Qj+hsrOX1bywS/sJORH2fisFmGG79anGmX8H2uhylWyFgH8b0LT1AoCi
HM3gbRDNeDPHfTUBoOzkPURpW0KDn+a2Wu/gTkRa3txsnh5fGNuOxiAPIMBAigkQbdwFMui7anee
SwoF91+9gzD4p2cps0WmIjnb0lbfAPHCBScoz+V8s7DzAGlnfLwfP8pJaP9DEPXaLqbuFFWxHtft
DSje2YahWeGSvdpE7FLia328vIV/Rc68Quge/PWUQSvYwHAWTs27UvWBEtBeCL5vKgq/v127uOg5
hmEzvwNNP2E3htK7TZGNHkrPIcmPz1RUBzvCen+vaS8cX73zzr1z++ew6mK7BuioCm2naP5VDlzA
x6b20rv28zwDbf9+KsYjRGUwD46cH5Blw33ymZ6WswmR9Dtil2LVHli4w3m34LnCIX7N2BMEGxUG
fn5MNs8UksDN6LxmdybZ90yIS1UVS/Qoy0dFgSzmt/Q8H8ug6XKXdcJfyZaQKqZSsfQVCe9KgB2w
we7ACCe3f1F/L8b240axEDrvHVCqpGPzZbzLmB4d0bBUmFyfRHXICOdIy/BGULlfXxTrOGgdAb0v
wO8BLx8FuMjyvDNuO0MrFVph47ioABUIHQ9YB7QlphrXmPKaem8abSJfqmO4qAelz38rz5p0zTNo
dEY7aBynjsahOjPrX8SuL9GDIqEoqLtNlNUfvVNRVOJmgkiYxoKET4pCvE8gZsIRVVCJTo07ea9Y
QdPgV/UVkogx2cLS0HuYNKzu8JxeOOfWYIpfxI+JGmHibHkANuZUVbNrMWwu/v0VHL0H+L4r5pZ6
eMeaMXpjC8fhLvsax/jBJZ774DCl23l4i6I/KN8DNloY2IVTyspu8Y2+xE2xAAnwo8SPc80JU4F1
spAworQ3T5yEuLg++drby6A3Fr/5UBQ0gGpjHAH53x1ZBv9ZAovAcXhOmGAsGba7OwgVJhhSs6d3
84xktMoenbjE5m2l2CvcmSoX6YGQB2z8w2KSLBhizjC10zmv61IySNGJmxyCnvvT1FFqExf2QLow
eOQ4PPqhYc6FgCK/sI5cerablDig+O9yOVyhRXKZXBhdyFnB1do9wFjHs5oeuPLoKZTaVTeNaEnt
tKX314CRQ5RvJDON12oJy5grCiQsKzJXP1PFEYrfIvkOPUvH5+kZHUocf95KiZa9k3UtWR1wPnuQ
NCvCJtzCLS8zU+gdlBQEIlPSx22tM2KAJsBOuWRVkVHLE86RLMBE6gagrXTMuSSxmMhmBqHGanb5
NN1YZgMUHMrlHLMQdQSGNA4z97Q/aaGQgRhNPU2vzrXDu5uMeCO735wmaxMi1jtWKerw7fGSBG1P
CQXNPhjJve56X2UtWTitG1c0noxzF5NTPPxGv1WL2lOwe8vokGPV9O2IISKkyCRw4NKI1U/JFv0U
XRyMVMKvFP1AZo502rUSbr4doz3m0szqY8MxAe/9G1s/Yd7WqUIbMi+VAembmjLmO89+UCQQsdDB
EiTQZU192VWQwtjEhz/1/O+SrZiN1p3dCKRIVzO3FNie+PofWdbLd2JNgCG0uTYHCt3SiYXbYxfr
y2iJuouiMuz++8reetNhyhjdnXVKE0mFwcO4QVG6YDIymRSZH5AO6cyggSiOzca4TB8dfvghMKFp
zmsOJ5XXkrkPqWcnYl/M4LUV8///hpRnLornCGmBj3wHRs3DRLiJrzb8deNxzEVipBXX8JKcJ8kD
ZtuL8crsL0El/xCxTDXmb9ygSbKBr8u030OtvrpXw9wKQmEIhHst2VZENMgW6EEZlCfNh935CVBV
6K++Tr6+fAfGZqiKfbMCTn0UCwMaByC90qzpXmBgwuQD+XYyfAGHFBtd8MDWSjAMafY8/ALBCTBj
I/+U5zZHVsarKqD8njJE14zQzDYlp1S1rQ+LSYFxyo/3QGOgj07JuZvnYzRRfTxdYN+ITcXBpz3g
bGhEh6TSH/eTkN8mLcFALBKOXmBSh3+9WyaJuM9xbNajhLwYtEGFPFSl0bs+RQa21FSFHzDCR1e9
3uyoM6MnmZgubg/sUHvRkms79RVe6wMKiJ6C3gmjrtEMMVey515E4LQ8QUOmV2SYtgvmKA/RwGoh
xk8iqp1QL6oCaI9U7nlgeAd1kDDDqX1Doy9EmT5sh5pWWrChP88Qm0AbwR0TOoVGkEMJ6rJ8ia6G
yX43wteTO8STuFClxHrq68Mqxol3o5xGmGZjWXpRTMjbTfcECHPDuU+r7LVQEGzochCUBOBTCy0e
ZlouOEtamJVE1gE7QQO6bhJz1j6zZuePITsOX/jfte7S0MV34yzo2aHhO9gC/cNYTackDWeXHIu+
48KNIrkh+flIhuEYfdM1Xi6TUZIQR/ALJvuGSJVpNlpsp1AhTDeAdy0pEIhx3f1MV9xD0vCShelo
4R60xGESYB2te2qG/EMSWgmBgOCE+xJgsVggvwanxAY0CrDYsXY948DBUzAXjodMmvm/lDCDS1hP
crqftRN7GAoIBxXGpWwmr7r6OR+0zRozsC2kYcTrSNuwDTKyB3aAiOT4UbWcR2MGIrDmdX6QaIUq
gMRYn6AjUEKfI8D2NPGmwlKqDRydjyRQLJbFoOMPP2fINmG+cK3qt/rVOSVegah7KF9wzuw+FA2z
8JHOywEMtVXjS36wnt0MnUs9JeAMeHfimqtuI3eBvQZoI1ZrbPSCkfYsAovFB9kEguNVz4Nsmsvv
IDh5E6DfqIOiNuosUWCbO/IbG8F1mMBfCSb4eKq8oWHLkrcMXgZUeO8qzVSIbK4vbg4uKlqB9KmM
8MUh5d3+SXvNn4oR3eiFm04Q9w/mpm4jWJri3TbEGrCsEuccv3rxQ+qX6YgDLoKO7LoHqevocyqY
NJt6bDy/zpEtT3w0gDzz8plQeEAp62yB2U/Dezyg/vJsct53KgN3VVORr3+Xl1o0Di20O/CWpzeB
3k49dpHa7KR9B/H76KdJ/k2QOy8598wDm+TTfA6ftaGS/OPdrgIcl1k6ip4LV4txtMhQo15hRUXx
OgMdqSXwei/zMuqeQP1NOs6zmlhYpAuOAxFJ+BFG3FVugL3NL5agUnklnQF7GebdgQ3ZxcGvdnk7
04jVh2672Pkbvf6A3z8NHdf4CdJF1ypDQ9XLX1zMKVy0NH4q1bAiJAGn0y2gDCHyWnu+0anUxn5P
JX+Z7V4cNvcV2ui/7/k0hGC6kh+Inn+OxXDZEU4q/d8iVD8PxO8rhVk1SBaRqopBP3xoTy8w04+n
xEACrlkZjlJOVL97ss1HyovXTepkOtMg/WV3BC/3c3f7nWtUnoH5zUQmWMf254IDNbdn4abtHx2b
5KhIFKym5Lx8bAM9iqUigwbJrDdubkbQc8Kj28qjhRUzyNhLNXc6XWFVowdbtAf8V1ofUauuvFZr
3DgpUrTOR6MGEn2fSOCjedEbzy6xP9PIolxWWIrk2fCVMCHNzZNpbCfvBn3JsfLCDDQ5lhDtfNra
ms+F+UozxeuM2rIjqahGSlBsCnRFL2AruC9yOv5LJdE2Zyvk3T4WTeoVUvg5sB/8i5g2OkZytC3O
/UfF+yW295ms68kOZsximxvTvFZIB+J8N2uyXTvZ0BAoGqjr1v5g1CxA7flIeQv1AGzsLBhyy/cO
n39zEmZedYok6z98R6hEVjWzIem9sKRZeOa81UinYPeUC47p9JeoYraJoyUSvXJJoBc64CQdqpMF
JhMwjCC1dqFxXGDOLB3wmfQq6PNjQqVHMwi+dYzxFvnjsZtGdEtgaa6KIDfKfc+jKN1NC4ZMjti3
fDmp+lzkmhgELK3el2y/vQKpt3j7gVi6hiV+B2p5fzNQt6OE2F2VKMJl23ch/M3bJ4/NcCRmtooq
7JI1Oa7kaLXrvQM/wdR/KSJ74/wP3G4d+gsrUWeZz9/7mGl0bcRm4YaORDJm6Q8Nn8j/qre1FPRM
yYoYg0rJpAhCvNPPtMfCCLuqNOrLuxK98lXXyV1lGSfwunTDhOdP9K3Tr6QacxqRTTQ6qhXfFRy8
t9oBvuzrNIFF6QVLS1ehLdmAHfPZQUdbPavAyvr04BODQUsT1N4VIOjb0QcPYoUrPBRXn7r4HYBe
7B+jAAjFoPDSwqBB6/jbQK39KkJx2LwWQNpzfWy8lOTXbd4MV7Tn5osACAGeFPAB4ehU8qyCXfqq
zbUpUdeOlYdDY+RmcEn4Hkjeis8MF93xdlVr8X3GZcTOqMgZvNL7cynI8u577azAprIiwVpUR6sg
oJpRNDbXXOBIgPCcbWjGudZfAdnTQQmrS0tbKwejRyuOK/29NrzSS0Y45yl6oESRrzRvuxbDKuD3
KweAsUasaqesg4qu/ksqIRyLPgZeYXbF2iB3FqI30a06E9LxI80Ltud8E9wbE/cvFLEKxAJRlpG8
yq3wYsIBzTaS7xEw3bfuQE7vPkR45ocfFAZVyH2xWyrqRjd1qnolcWOqaNzmffVVthLjfOx2Agst
VGxnqXyvxj1pmnMvEdBzKG4rtFGbQI2mnQmEtSc25DQwErQwmhceqmpdPGYEsAUT26p7TknKzJZm
+C5Up7eFX39B640HzU6fXHxwQsv7yjn6GZVwpvIf3kMPAERjtC3M7PLwNMcirvWGHh7UV2qLTNQT
gIlizn+3nM7YDuS9m2wZmk6M6zDCX3eyl3f40sHwoqiQh9iDmf57+HmWoFA1W+BiqRXToaybaTu0
aa243KIAxRjtxyunBaDfQpTk17ldmKSMPVUdeoLNIno7jTmLbEwJap3j2KzBNBHi04kaVUIVaonh
3u30aNKUlvelMZRjnUUy/CUIagbcutREhjhpPyFs5l5z+VCZca0823BzafeRuYXo7cQxkl2Ot6Eo
kj+skKQT17DHGPfvlwUiM/KXcmRJz0P7sLKuk6Y1JN7SrrQlv0MxDKE8AirmbpkfHaaNS4q2tFEE
8iVXO+g9m8q7d4ZHkxpjU1o0auyrGqs3+D7uNjDI7fr/1ryQCLYS/ipgzymeeC1EKy+IGFcB/h91
IiOdHzrn+5kqG66BgVSGUfieXV1MjwEWEvObVgwltXuLPDpnX+BHt8zB3gZQXFHDkkWekbSw6U02
VJ3hzy2zw6zRChilE3SgVyybLQ0Wp2zS9AXYOeN23Tb5FPFDx46wMBpcN6C1cEC355kNZFw7vGNk
HUlxqrCujxQDLv4hn5MJ70yqDQ38j3zLZZ15ReYqAtIE5lCymlMhVHVx+VZWqsuMYxg7CrQasIKO
mJZbOpzXoYfeThcIqDvZe3fkeCbhGePFUuSAzDDcoC3WUxB8Ge5Qr0Quwv0f5SlZ4p4w6fYqXqPR
8cFPRpfiQo2goMKESk42XsgTj5qalQGQE/AhYA213Odf6SxA2X1MQtwwldjXDhXplrj/J6Q0QttA
7ir9qqKJcvyNdK5URhE5KXHrk3QYBMgYJeR+eC+ZV0/H58Cx0Bp2Ujjizv4cpFrpAqAcDQOQfYsl
OWcRaLFDj3hT4QfAoVujxa68AHjS0Z57BFKwA0B2N0y801uM+yamS8p8Z++RQGffykbBAhVvM0FY
3jSrhvUVn5J54Q33J9UE9jm4AntBwikd5541y4LiQRQyF9KtEm57gLB54YXe9GENi79MDOCqFCrN
0new0wnu8VMIXzjFf8SjI6Ntn5cTt9gNmYd9HFrQok4z25TbxUsip73MYgXGLKX8R53VkdnJX5wK
uQn7TCi6KybjVrJMEKNywP5L9i2cjOWw2TEZzD2ZnWrSTPQF3jkG87fGxJXmgPvjRp1uVAQJdDPF
E4I7FrAiXMg92Pdiu1nsOlbYKl07Ljt7CIL80R2xAcQA9/X3tTgW83sT5jnejN2HKoq6oyCvbAdW
S6V031nJodLGkIXK5ovQUnDOpSbWKQtR3hb5gYiRZfD9epjxqw9b/Qsnv77BfVms8Mx6SHHDDruq
U6p3X3nWx2Tk4AkF170RST//DrpxNlI+2NurK1tFJ9bUH6qfvTO5N2gC3h8wJWb6NEvPuuarPfxa
id38gvTVhTKIrY65CbpOx6DGlfiP0RB3cLHz6pVnTZf586HwT6JcRasVVO0OmkWbOsNLdke6XY+w
rumQpIw6Nz0hvKJek36oyfhDcZFuqL2Yk9CpkjYf+5ZX6/AKchwMfnlK6OFnywCRlmY4yx/TqVdZ
vWwufwW6w79QrSfRpW8SAG7uon5USCttITVFa4p36V32hb1kjOl9OYrQy8kPVPV7kudp9446zRHN
+EquxIODida9TOtdahRFBEefD8X2huUDRuwqVo1Gnc1eCnBmc7KsnvymbJF0bXc6KrlNfgk4nmuj
iu+72ZHm0Wqf76J0+8oBhiJVZzDCmZPvvGsrCx4quKvaozlSN60YSmXAhEic6Asv7Dz3xLq4PZNM
3DhAydP+IOhUc1uXBtkOs4qUW8U/Q6t8TsuddBYRi6FbqA4FcCd6giRi/2tKKUjMvrYbvel6Qn7U
QaQs/xLGY2e67qLFkSJcvf5YOudDz4RPtLrMzAbkCSFe8OMN/8sJHhSw7FdpvQ2ZE6gJbh3Sr/wc
aTdw7g7sahsP214LwlTybxhoo1JYGC07BJuptnjcb7DSrWYh84+XC+xPnK0gbD/FPHRjBZ+7eBAS
lZqYKGtanptqw5yXfOK3K0DXl49pME7BQsoF0IixYsBADWxIJsKQf65Jtjl08SPYFPnmkhgE+YS5
axGJbl3aGF7VvBSh14mdxaNvx1iHG0c1yMB7PztYxMo5U22WZj2kpJxXdaqPTQbkfhUdGHWwSi6j
vmjnPptiUB/qw8UgpDU+tBTX8suCuWXjT5uvXn0MtUInglTHNgVTA5l8bysbBTepfNH3hBOk49p4
rv2L9OU01AAE0y4Lb9Goym/ODkljbMc+cPtf1biN/ytwgPgHVF6Ieo/pVOhaMzTsmbsoUbC1e00y
FDPCq/74dsWP8dMj1xAb5YhEPYsoO4ckKxYUS2/2CV8ACDtnUD2wFrEZ1T4Leaii+HbwcF4CKqke
YDwC8ENQanSzotWiTbjDYfScPSvEsmp016Wn/gI4UbMogbWBQq3YoTLAyAPLo98zIYeH53NzuUlO
ztqbegTecuEFDMjSHXr6AGcXqrUlLx/iVvh9bAabZvp1IHEl+b2On12JWuOa+YmzLlqN73rxD0Va
lS/noim0CuGihd5eBwZ7JYk5Hi9XNwh41uanDiZxJnb1h0xq47oQaAxSg+Cga8V29RYvWpgTdey1
Wi4zsSo8J5gjEooW2Aq2WBdLsNqcYmrrFqmGFe7AIrjhkC8FurAcb3LnJG6shu8q2Yi1198w8IfL
Hm8UC8Q7jNgaSYylLpmhsIz10NyyhOiOhLuCKEdh/aUmYS+fe5a0XsgJrNt3D+O823f+T1+VzKG3
621+hKkz09Ia62jGQfnI8C/dXi/ijr/5TLiCZQLB07oklk9AnA3zaBTsyRFjFH5/aKwu8Q8whxoG
c46YNTOm857x19UeXDNnsLX4dsSg/TiNYx8NNHUesyt5mwUET3BMmSfiBAki/vDrDHqxiO+V5oWN
kxvAg0kNS/ZFQMeFkK7PV7wSD9mr7UjgEameOYt4FvSMsJf9vDee3/5S6DBoJf6e7crbTzeBX2KD
sPgzA7ZxFcy3sLBefNMCcHHE7DaA+GX1MnKANUcvMR4gLbg4neNJptaUNaaq++0iAndgJZMmav2L
dTDg4kdHNV529iNq1G0hv9tho9P1v24MFFju/6lYUMNlLsfrRieQyCZ7s6JAXKME1qfvkwa7B0CJ
aDxNyDzXfH0o94xVyfeJ8ZWTS92vUx57U7t2gjDyCGmXCmh/5ZlIqqwQA65Ll1GyRhhAVShZpmyD
dmIDC080LTQzpdc7KsKxdAbjkAU8cdAGip5CHZVzU9cwC4TcpMXm6FZRnKDvTz8ROKVqlemZ/PWT
wtQafwkY0xRzj6/e3S2ELK7wgsucULS2AklJzTHFTcOlaBKHoQd1+Gbnz5nsOrbUEPApI1XB0+4y
tzMMh1v4OIl6Sk/0R0Ll8Bm8H1NSMUSETUS4v3q/J15TR7S14NbeTrSbAYtzoL2ivP1tWkmUQR0/
fA3C5sAwDz9dcG5t+rAXQiaxTgA+O54jHiJzX/hqSrNZo99Ddi6g5Z+ji5xXNwMdNRculcMKg5Ba
cgxKZM2bhjNoC57mXIiR3frZFhFg044X0cxcHBUbrWPx/5uMVgRZV9Bx8xE4+tTqq9SOoYtN14oh
DlUqDLE8YAVoniNprj6LxIv+AMNenjYuWP62nyv1lb4Yhlw6f04D6IdSzHM5euxTjw6yPgenW8c4
cBvcORDa7j5czqcF/TP9G37onNpkbaKTEvy4OZqhpEtpc6fAgF/rivxJgZtLCLCRfGeNX9wDfr/0
WQ4TNwiusHB00TD2Szy9BtAFe+b0B4YBQJ1JrG7xNzd+BoNy2h2TXUxT4MwEZEEEvYySynWHpDmQ
HeGIty9TSDF01TkQgR0hB3kSu1XmHUulX0Abf9JjJQn3xWx0eK6co8dKyE6IJJGb85oO1sfObpMN
mG+weQvydHvU5c7Q2EI4gBZkxKBnBZWZ+eDb/XIG8m82DSRKuaeFCj0tvXnHqyu6LNGPS5KVZb+U
yTkqWdQnePcWBMR3Ci3YrvSLC656SyoM6vTVdwXtI6w1vLxEkSxXPObVzgBP+VNuhjuBDC9WwMzz
J4VmRisXUsZBFV+0YvzXKnM7t2dDdUPNLKGthlLI1lAORqE1kpGI6ImbSH0XewXsp+AdMLOr6GwW
IdfG7CghpDBrPBT0VMHAkta3Vd71NTQtwqnHeqSJf0045UXFg8cL6IweLA03VCL1sNJS2UU7Ue/T
5NaJh+vuR32jhiB3JrgVksMvg9KvVYiuENY8wCbf6DQOODvmaIzt19jD3zbDdqa41XMlr2fE21xX
0ezt2b8Zb9pwBQ3Lufswx3g/kZKP3iSkYiq9voiAKYo5BchyQKRCa076Me5rU4vpnqvy0GiVBCik
3dUnShn6XSmbL8lUbI5rA0ySYBUuSB/pufmgegAJHqOsX2tA9/SGUVmQxUwnLcFW0pXK7MoZnojF
w5Efi0OFP9omDRys6391PyWGUGxkB9UZsIU88xboTTpA5DHHyYi9ALqgKB0Dcgalynp0jXiX7Ycz
h/06fj+1z07DKUNrFQMBQV/gv0gsvPJp3zGCySogMV/D/U+SpZM9m/GMzyyqWdKS+gVMV2UJjJo4
kO4SbA+pLkPEYqF9mtXD2FJyhgCSgdyYSQd3pVwaO64tbD6s6qs14WYqhP2enrFfHCr5gKQ9/PFm
J6jmDUflx+Xo7vtR44DUlFmEXUypgerEiSl+L0dVUSFoZd19f1HsEKSVH0QUJsxnsnTjVnJT+PNO
adhzW+QqEQACf8x/kYtLMBkcpy0OwyafSnIftgciamz+UVVQ9BXKH47qYyOQLi81pCErkXG799wt
HrNYjJ+5dDMHYQkL2BXfYBsYN7ecL5JH9l/ip/hq9LS7uVEdw2PXV6Kxn70xRWOUvEzLoNiUSQkr
CVWJidAjCaDengRuZixRtU/L689ACiHU4qZhBH3p7HX+SPvhYX575kngWS+ukifNZA19Fi9/eXyL
5OyLRZmkRCg/rylty1VNlj7pjMRrUpCTnFmcMGXy0LMqeo9Twy8eqQ5lixgOJTksELW29OVmElGw
kcr3tokZ6IjyvO7aaR4wio4r0xvJML52dyQsAb/CIZQRumnDcIZu9IIgRRhAYeq8ypxXRMk5M04U
6g+cXOKtewWrCQyV5TtQqdasOjyGYMl9yG5eZxPIe+uLWjCEVoOLhbcZoLSjiwkFKP+bcVZE7Hd2
VvxtAEDBqE6Drvjx8eMDSdOqAPzxGGgeMw4nsqzIbC0UabZ6CLw44eXj2XQIKDVLxT+Vz4GNpBW/
l4lH6XRskxpJIpYTB3O3uhC5OuMJQfuF528LMvqTb06HWKDHCR54V+1xo0G3QbSmPJOOWvVuZlpo
HLhsgjvOBiz+q/2zNP7uPWyOqV0nE9Zvy5Fs5R/Mh4qkQoudha0d1zab43hTFK53Q+k6VYBxKvIe
K4RyhFEAbVQG+4FKsCBW3JiUddazhyFUV0faa/w8PXW6dGEdOhdydu30I/hw6+b1Xq35aBqiuCSm
7QmhYvSqf+S/Op1ffw9KU5LLfBbvZr5nMLUro9CSm4qtPRqJAYKF3Zm8Wob49Air30wj3bgRZDai
hoEaz3FF4opTWJDg0ZP58TplD9RmThAVrQdoos29XmNTkWEZNksl2mPpINW5ZHTKPDkolrY0hsUD
UX2Sbd+2jSPBW9mLyeVWDkziksx39wQQmcfwe6KPEgrReC+hHfK+WUEnZu7exUyC9eSfvzKiFlPT
lPq6zk7F6HXMIt/ipZCB4hPWwSq3Iy9iIFd1zT7di9JX9MA6BB70BanaEx5GeYQXYfHnG+Ep+uu1
UpV/K1f5gZEeyfsbV0oJRookWVQIIR5QTXkvsC3LJhNd5QfnUu5hQ8XjotwoWWo8JuNzIFcTDvM3
OCOEpwuqTfjyuDbisIrXp/exSnGhyporPzRFBDGYa5YePrTjEoZ1Jc1CwUcMKNYEpwl9/gEXBXfp
ZwXeb7V1nJ8gNJ9satoISpJhRcqEYx1lD7vWzAinOJ13cBTB7MgUZcAwcLqiqH4Fs3je4O901QuN
PjPIfbDrKL/d3HMWbyt8LCQtpldtsNgx+ORiWsSNZeW8HZbmbMyA18KVaKz8aH9g2mll+Bn0oJ1c
4cQ474T5wHGtfH5kGvZl50lV1l5HbaxFSZ3KbOCBTjr3A+zyu5QKZvMdXKnkv8b+XS+WHurGNp6T
c0gpaBbdrRE+27DnJN59JTRuXmarUO19Z+TeDWaZs1qgigmeQGT+2gc/OjhNZionLxBDURaoIePJ
9/8p2nII2DShULyOIqfvxjpgx3vcCno3rE/1uKfu1Nizu6VtFJtDLWaSyNKhjG0jjvgkuCvgt7xR
t8q227bL5fvbUAlvnn3eDJxx1fEiKc6Y3dzQ3GgKX69qcmrfkJjopX+gqE737XzWntWfrgCDh+yC
8Gh1UtjlHlw7CVn9xUyiPyqJRk075XPME+tUGTZ+A+i07MBgdYCXfMHfYwkt5mS/preNFgzPBpW/
zM6FRQBFUH8ppHZjSStYF9+Lv/ZbsHuHKzmid2wZV9LXEtLjtJXDiqhJ3L4u/yt9D7GRtPdkiRYj
ZbqxlOk1xohQGc0URIMBg90nr04zA7mlfDyjB60IgHvN6H0ih57MnHl/w7QD9LrZuPAXW4rnT3ub
y+1BJW6GdYI16a2njnfjQQld2e3tYd8nZ9ciQwHNW5bnftz5DhF+zATAg42xgE4OGFSY8iJ5qSP7
wgy7QkglwCSgpYflJ1VgxGRJL4+Fc8wNXrhM72l3C80LkfhrvVio+HNg+qBHhNs45rcVaWMLs/uh
iHOueRSJ3JENlauvA+vIKSy/kHYnsbCUtEf6qx/NSYP3q4RQ91uJmInVRMS9Re3GOJbwZiyXohAl
GTc+CSpx4wdC8mEUELG5XXM8/KAgzBSXdaQ++JmCgCrMFrnxohAxftXdWjx5wBCqdKQY9zcim9VP
5tCRWhWUDHp39mDXOECEhKBK/uslc/PB5lou7gtNYXHFR6dcotmb/liLwj5N77lko2dMi/zwkSzF
LErT2uf5kpvOWEKEqqbmG6A5sD9D91jQKNY9XjPa+bx2H/RsXQIeFPa9dKicfW2xyI8Svfq+AOxe
jTF/aJuqNsUc7wLHRPyIibJwUaHbT9eIPdU9oOBvVo8SY3JcvKP+PX1GBJdz8W628aLKvyNYP1U5
6s8/PJpOUr75UFUH5dxArtz6Vu5JWPRQvRBcg35eAlD9JjHrZsrLqsEq4Qjju+M95BMOT81xxCgS
PBaN5gNKsJNoCtWxE8ke2ZDMw6Ro9c3k3VB/4di5BpgRocbIK9XVOSt7v92RhGyj1G6s5+rb9Sw9
5386YuHZgYNzHqxGUku5OZfUWMprKhrxnHZ7kSPoSSwN1ndy61hZu3VJULYf31siRcM3Ohbg8+um
oKBODkaVh4CbeFc/bVGpoFYY0XqRvUt+eLHhXBZu8hU8WEaU1OFYGKOxUZ2mty01YiRQot+olNXQ
aStiJ9Qqi+rKJrZ4bFt75Nl3hacCHw9GPHb29eTuf6gmQk7bNuJ5zND8MFnzw4x7WD5PQ8nVXLaK
NVPtjOO+UDpPwmGcppROJGIelyW9e6GN7f54g5XDXABieRx63/ViJCW94m6+BvYk/BDrj8wmvC9g
8KyMggO5Mxbi532b+hFP+/dvXS2Vm6ZKAwYvHrFspDZYJ9aZU4hctODVf5FkQaULGgIJU4yx+x6U
AoVBpXcY7bUMDHOXjDOe/q9bu1iga3lXWm5eDBE8aWiYP4rRHAefp/eIoqSj5GcxPGT1r/kGkYbG
5qe9CA7168F/lcJFU94oiZpNfpWPCfjqbKR3F+yxSKz9b/a7XSaDXp8kVaTdzxFzHWEjJb2WytFU
d09pbEdhFca2Fypbt+O208neeDlYwxABtr6wDDntbZa/hTou75kKqKLWLBpyw4Ejxv4woekLfTcV
1fG7/NDNpSqZY9vGX4iKAVFx6eZ4GfBX6PgtgTu9tdaTXwEDM7Ya8Ien6EER8WjdjfEID16pGsNa
Tn5FFQR767UmhWMj414lzFeX+POjswLg9ClS5JvMQEIsZQkF4h/4Ct4qOj4Jfkn4AKEhsfBi4Ypk
42k9tm05HPhABH8R9gvWOcpVKYJLc5fZ0eu7yO/dWw64r9Xt7f7zQiXYixc4pK96CfALUmrAzRU5
GsFWFFNB4O/3gmv7/ISfLMR1hJ1eOeYAOkZrTOwmPQUjeTo9rI4c1xKE5qWvEH5B/besHmbGRqB9
IVQqP2izBtSADJP4R/yDktJbm9zw5WkT/sZIcyRQWXObcCbEORhop4A/VNDB8O0oBbcSA9/GEBnT
krWSkiT7Nn4P+H5liceM182yyWvnu3da+kFgQmCfEKpkuMvcG+bDO+5WWoLBXFolqGzRxQYWKqHb
344DyU6p6BZ5aoCM8LWvdQADhcu+GV6kPqlml+PAUuoxOl9jfD7Hzfk4A5GGbyPeTnO5WY7tT9OQ
vxCA/YKmyq2CB+gbzcPGJTSbLF3hg7P36AzhXk8k4obXkD/RxwhhOmIFBm2/vWcbze5EvfOYpiVZ
swMIZBEiKy4lOHDcq6HBpNRNazjheGLszbNzaEXcNZHrHK86M5ce3H8Q/v/p9cETTaSEM5+XT8zm
R95SJ8OwDWTmsmi1kHuD2x3J0W4M2swq4jx85yi2evFK8t2R791kdkisy8bse0/+YZOl32H0HQoW
bOGljZuc7Wg0XsCHPXBgQzvtWCW6mL4Qk93jcQOBYeX8GtEXy2roXb/TbFMt1e23vB7ZU8wuL9nB
q3/IoOtCfdSe7vJzuaoBYKAutIcDCEOAfZvGNQUgegk3aeANLtqCl2XeXnHZKAEFVwJnBZnNiP6n
qJc4PQ0L/DfakSUCA/f59PgrK9jveSHOCgaB93Dk6hhYNWCnCV/GX0tAbp2OlRPBoW9tRY1ArRhO
iSFoQsFQIc7esXjf97usS8LMlcCqExHJ4JRmHdEcaJZVvPJZx2CoNI9/gMqskp4DCqm5o95IDCKd
YGPUETEBiXk45scNcnbCtkSYAL21hrRXPFtg1kCLsV8ncfmZ/OI0NKxeJcifWZdLtRYieNI72GwJ
qlDZu/7rJKh5F+Ut0rmfrrvmirqhflyVZufLx++m4kGc7rTmOQavBcWH7Zp4tPZx3F7C/RiGqIcr
42VbVQvP8KG7iVOV+tMVWNhPmQL/nn2bV4+biCUtsguow4HLPd2sTUs0LwUq1XzPEoVs6u3ASn9/
ErUrVnu5Smz5RprM3kq8kJLVRrH0FYV3iSrE6/F88Wd4mDiMsfnLwhE6ATDsmz50lodQUBvGALME
H8eGLyBI+Y712zUAQsbJQiQ0n3crSzbYYb6/AAyQvDwmQYORTO91XPRCkww1YFYglUfFtOlk3MMX
aN/zt2kXEJe4m84I8csetC5UpdlNadeLJubac+aD/tIesDlC3+hwU92xvPnx+bQnC1ibuN+0ZsJ0
eDu/0HamGUd/9VSgH62pV2vT2+38H3zdDA90/r+3CAwdgwnzDqbh+3WRvMrIgQ50eS+D+O23pGGy
KsP6RmKEQp1riS3Y6V9gnSEAnVhRL1AUSToOj4AvwpzRqBdqqJJmxFuXre8w7AJtu52MkO5DU25Z
Uc6nnI38qbc/0bbcCKKuxcm0cJ/MT+OP7y5F14hr2okW9FTlG9jwxKXhvVgP7t3gWYeGuTk29GR0
226AzH0Cp1lfENzNUplv5E+lDbFS7zlLFWwUzbqfvH7JsMwzDc8U2/FEDmZJahl5ZOM/EtaYUhkq
C3mkpmRWEjOsCrvY5Gpyom8JZFAfmyUZFrtD3Gnh8ng2IewCTq3MNRUM3biSWtEmtu7R8yFZ2C+n
ypHJG/H5DUror6gHhkujvvuJH5X7dlJexjXmRvzhyUvlVz/o6vNRymewokVwUbLBQqCvkHGhdKNK
ynV1SfOlgY+yi8ezWUK5JYnYEEUC9i8NXa1qpKVjXydxeb9OSQa77l6PK6ghPGaacx3be67zkTJs
2XSkgrQLx5CQyjy1r5J/UDkONx2FLEAnWLGuYMrtyZ4DpelnvRT/khherMvIzeM5/ggVfL73I5mv
8BuWmfr/gySlD5ji0yIOCaXhDRAMVJP5sMjDtzwq7vltdnlwIjx9h/6EsdJa2Lh8CSBmH7N/eCHP
1jcfYmOiH8z6tluL0NCHXAqhOHA6OVpBP2mQD2DWs2ab/dPX0XR1zzrH/G1Q1+o1kwwMrjIj/evr
rVKDbSuukQ1p4seCEoVZF0kKncOwunpZHyf9GoBaXDwhV8zkoQwWbXSwYmcBzdhQtUFMkd2/AMoR
Bn0Lys5Jjtyj+9LJ0BqElnNoYejtqDzKw3qC7m5d9JpEB0m+DCR+dfT3/jbSuMvtk4LSH9MPq4C/
Rydu0uO9ZnUy5rSWTqBTAN+v/sfXf3FarkPEezwmp4GFI9XajY9P9KXqBAb7V2mTY/Q1i3h4RUpG
euQAwmH885kG4lxm2vVarkfA7X11Qif/Gi3liOHK+kFqvp4f8/y/JcUrVezmFp9qGwXDbC20yNLi
A0pf/hhvP92AdlvngEftvCZT6oly5sI/UMnxo+COwtWiTUBrYQ2hVf1bBb95Kqcvpz4chve/t22h
3DR7F2zg3ShcIei44CGZCs3ymGD0/F5xz7lsDL4fF/sypCU4dhIOOvYy/SETpZY4laSx+NVNYI9P
sojIxJAA/uMCr+y2Mi6xPwmuaYwzMIe58Car5IAdVMrv1lHqvQBBFgErUV1B1ihMyzzyu4F4pArJ
5+V0/5XANY2YfDVbptJPQrlYDTgn01u9/UVn2hn36SLysONiO/3YXnTMfTKZTp8DpBJRhoGiSReu
X1E9WJPl2WR/kIoCBEfrbpqmTVrrViiWiToj81NgWVVDn8s3w9nKFjTii1Gaa4Bo9XksrG+cGVsA
VWkTbEm8343NGD4x6eTNr+NEJSdAfeqmzTS72kLbPrHucrnLusv6tLpAlMjMwGBcre2mwCwYYMOU
6PabB6K2VfdHwKDD/f2jOY3iyUW2YkOeLQSW360/bQN+F1lkcVok8/eRnT14Mq+bO1f4l3Re59U9
Rsp/KITzZ8mBcqWitjDDIiYzRBmtOFDFtX1PaKBigJtVX/7Uw3Blp943uHrhJ58f7qaC5JnA3dmY
19aGGAjFD4FfsYqvavJUA6UYdpWtUqAKz2o85hhcICs3JYENxeur+cPeJ74l/TRkBRbRIPT81Q8z
sgsORKrFwTxyEfYTtRpjvrVOE5igN0/MtJpM5RKwapRjP6WAIKaVIcc095yPY+0EvNUQoMjtjG7z
xX4yGY6rWqU27Rz0B8s4p/GdN8I9cOOj8JDtjV+9fx0QZqaPa4PgTN7je6dr1UIU/Gd7InY78luS
D18I5hmHOEpay4j0h7HEDvFI6focPU/cNGB8duy6Dvt2O9yrxppxege2lfKFf3Ryd9HtHD7Y4Q1a
NuhTOQwXMf8hKLuZ+Xq8hF2mprMitLyCh9OnRNsDRkHLZP19D667z3Xork1MFEQaioCdqNrPmw5v
cqs5JMy9mja4yn7mLJX5Oqxo0IKfbZLK0rxWu6RGOEEJsxwFyiqGpNDqqUno4BN5mo1V3e3hBf+h
tOP7ajzGo9z35j57P/hCOZj2uTQaroPm542UZ+SEqmMoNAAmBTiQi8TkkB6B/vTxW3/BS1KTv0V/
KHH36w1DrSamUY4Fa+9mvqte+XD+hYZT89M3/dKcFyCd++PB22d7F4MV5u2ZdkydZjgUg10GiEoG
shqvW/s+h0tHs54ls1nM7egu0HRlDhbxvPD7kbifLiPzKgCI5Nveph5y2nYcyoSA+7gw6ZWYvvWL
6DBWz3WfFGa+7960ikI4lzXIqADi3GZQSVR634qZgloi6nWODwWR4wNa1M3SyJhCtoIrKpx1KQhd
Wy+vAHmVPGPD+7O0ZfFVJ8lUqGyQTTpKGH4voD54yhFk2hBtOOi7mQubk0Ktox8wLQfGBYVQqUBz
1ElKt6W78vFdqTxn4Fc7l/CVaBrsaqURXsW17W/m1g1AmgGbDuVIoF740PjiZaMjTiH0hDerY/n6
8j8pNgVtblJL4/AbTN5itH13nInjAV0suI/NvOpwUMdHRmNgTt7pJDdc/VXtEygWfiIr7CIPEIR4
Idi5ZQxFyFJ4vU3xrByEQJCC5FKuVJ0+gCMWheXRdOQli2EHxjadZ8jRWFFAncYRU2LdLp60P1Oj
Iqv8gM2hhhQfM9fFliT+1ZAuQDAbLfkn6VEpU/3Utnye1NmJCgLLr4ksKfTGFt9Wvc/q+o4SHqGZ
qcXyp3+ToB6DbeOd/7HUB5GU5tHWA8lChzeq6ezhNkP8hPbgOiEsdl0KQLUJTYHUGLnuS2r+zGHc
YwzUjmg+d3fSwi6KSpLy6GlV3B5WTC8jew9SB97d2mVFBJNiAgMFGPoK53WmrnieMb0fVPiwjCFm
phoXpQb/UGqxrL7+gl4vW52oUmt+CuVLW8nr9/6ED0Hu6KnEs9eTIK3XWGBDFqIHHP26p9dn/fH3
jpoy3Or9Yf3G4rXKdkL2kJUv4ttZKSDmY6rvrfsf06YdTgPIbCQT9pgNt10ZoxEp7Xk9wZ9swz9s
jZa5pUex2VdNOfjFRPyYsDpAJG1i+v0drhFcC7XqJ2z7Q/3m/yv4xe2sodEDqfu68qG70CevPR80
EzpmyGA+f+s7WSNj4S5kaw7XzQwWe2wRnK/V0xmR0e/ssl/H71wZ8jTRDH7EIL+lCLYIqW/OPvts
UfCtpRc8HBgI4SOUsqEDvZGxWhUhT8Zz0WFQJgsjxZwZDBAlGfMtdpjrccf00SA0ldG80URu+oib
EhfPp6mpdhODKwWgeeS/ClRZk11YpRimtjQnXVcJCCM65Vsnkiy+udLOgedCX+qcmkGXHf3/NpaA
Gj0IgT2HIbeysEeTpXnKpDIjlESQ08P7cLOb/TR7xvLUmSJlGzs19vTIy0dbP76BYSSO84Uub2fX
mZQhALfnPd2L3FCxQgOelJQ0vNpeQSAbH+4s/JSxXxVpbquYqPD780ybnQLkIFnTQw95+LPbqfB0
Fvjinz14BArE/waAR4EdmgPtJb9p9wxUdMlytEk4BZc4p4oANElBFZDrqolYL96HRdEopeFKHXEg
fZJ3IMzsf44DWwgt1FAbgeKCpT+cAU5nDH356GzS2Vf4kQO2EKpDzqPxDA9SR/amimLwVWs3/aN0
4XVGC4bH1fes/NjXXtEq/rAw05F8fPq56v/MQrVGGSOr3QGvUGvtXxz1A1c/V+TDuuQQhNLTtWQV
qqF3JZtQQw0acl/fMR3IdJFPg5YMNKJuLXVxm373IOtdWloDVZh9G20XldnwuZcTbNL6mP+SRnW1
Q7MZQW2VqYEtYV50e3RhRkGk1JT4jclXPZY2AN4kvnrExuPpV8H68zWLmB7OrU4UBktOKwM8rzgt
a+PMUcH4ToVxPSgMKoDF3sZ2qzS01XEUfYM0UmidIZ8SxjXJ07w8G0oqDxQUaZqysaod0c8CjhMr
NVA4FhjvLq41j9VL8yGnDFuyRQV/obs4o/I0C1N3CDFH/aIgtKtYtR3OpneZph5co0Ps3oxRsUXQ
wJmEgyYrN6/t51dHEhHrT0Rp5ZILGpFGRJ3HxThZxc6qTY27GSsJ4YtMnOyN/AZx5TrFhRsISRxv
SHZvnrIAXgYuyhYt0Pcu8SDPaUEaGzyQccKcLibaV8yoTb3RFYEsdLsSpF0IL8lsUg7CLdYIelWL
itPLfXp1ls+g5eHxlDMCPmFDOBDpWk8YHH+ygU3usm1/daK4wz19b5JK1UnHtrmFmCkzdC/saNLZ
0jMn4m53whyacwy/m/iYxCg2zVvnhiWtoBWVdx6GC5d2N2hsS3f5zCnZI+7tHPacfneIuA22VGgx
NL/JJXUeeEuNQWMTnU1vj1ASSFlfGwFNqOyO/OYRmWVHFgfTnabcVf1wz7VXDfMjdO/NIjxtG5J+
1FzGAA+b/5aKv2nrDiW7jkonRRqVQT8sB6k7sSlKKbjlm0/0Qo8SxIhtmpOz2c3v+tmwqoTxE3SP
tOz9FJzfD4pKPyeIoo68A7VmuEA32S03mUQ7orczaw15K6kYYII1nV/L4Pr6JWHVhy4joN7LQxt6
UwnetK6gvuiTPLOCk1OrWKbl2t4Zu0ylupRDk73fK8xeBOdD68974uaX1X0goK9Wgxz5fqlhlaZU
VI92v27iDL/ENzwcyI2LuPbDT5VxP6vVCWr6F6X/tVsQnl43XmFHaGmy1SrlqhoOoec8/76k5vq3
Sno56WPFHvrVrDMYQ4quc+ogh8O7Sp6klzptb4u2ADrJfsNfVXbMzfEBVsWFrd2utPqAr9zE7B/a
0v93K27YqaET+XQEIAx4MTmRyq5lD+ZZ512doKjgw07BAULTiZ2BpPfPVuTiayClixRJSpRbHqVe
Q9GOqZK5GkdRJhnYlXyQKOYxwG/oaLAtpaIQhCBQF4td/OFtCQyUgeaeWp1DSuc49gBw7qTqYGkZ
Fv2iL4m+3WxAxr9BiHu4o3U8UtBrtkWxS0aBYkIrb9mfsaJTaxNBZYfXUkkuAZyRu9c0YEfqxmHh
UvPqdujCbGThPG5tWucNdu9aeBGfEeLfysjv06UiQWCs3UX5O13Rk03SaFF9s0WULxoi27O4YdJA
UIcGQS27nbG2bCOc+W4ZRWR5vV4GYHj+35oRde4uBqqVF96TQe2EZEOMOJcB9/Amldg8Eh00I4XO
Y/+dS1piWjNjTl99lHQ2yUl/VagIRpEzF2Ds+rrStlr/c9jqTEiPlTsQUbLHQPVzyOBVHEWH2/g+
AgaZFoojc84Hvu1Vtqfa9z7XlYmKTgJGfndGJKeAdP3z8UZestY78jvY+OZNdD8EGr68iueu3iM8
R3glXZqv+WEEYY3kkczcaQzI0QuZgDDm8cBoPkLwPPd/gQCHpDLeN/i5+fvfW54M8Pf29edSb4/Y
jgTZqyGGcV1MJ3sS7KpmwM23J3AT2d3Q0j0xJA+S7h0VRFGc9RP3fXwgH12q6hOw1ZitC66XAjBw
Gi4KscIHYb7W1eB7Go1uyjEjERjEY3gcSLnv7oHiKbKFNNB3CzizAjLwFdWsF3ImPBptezGA7FDa
eMy/4bIL8QRE4BRphP14hNq0wt6zI9E+XXevaG/ssdc3HUjymRXAMjHWY8D/iDlRSeTYnq7S7uQx
p4+BcteZfMWaE30uQ5JkeXjWzgHtyE/0toodsbHEPMLri7w6XVqeBfU2a0R1e3fGjCpAzNjeUjwK
CjM+TkQ6gKvHRGE5KoiV/ePSLVhRLEiZlBCqxNRTAD/Jcx2wMLzNlGZmNGsrg7tkHw5kzVZ/gGLU
75x3crkxjVnbET2nU2kkTWxIr9e+U0aiiPBeth+XNG/xVbFxSXhprb9dTaqs7356OTDuZsXkYUBA
39NWTZOEIJjc8m8gjnQ+fEliT74ceR3DqfXrPgitpHI7tGhjXfRnpMo95NGrh/4Yjh2tOgFxBFPu
3scsrFr8q0Z/3RfdlK9dObLP7n0PJFFnFtuWLQloYaqiCS9nq5jrJ7Efg7+5k1t47RGdINpzaJ/1
ehrv98k34v85XQ1oqAVxeeGfZG/9oXhyLl3nsfh/AqaQpyukJicyQf0MkWiuztK7plBC+sVIyxDd
n8JHnEZY+gAiYyCu92RSlbw9PxVeguDM7DPoI4AUBhGMaH2HHdztJER2VBGZvfdf0wBeBSAa2G5M
YAqXfIE9+mwPyZGY4wcu+eTRKQOvjETMis1xiM7TxOc584DWBLo5a7QSXhx8kKy76f8QMjKB/kbq
1m8fbGnqeVcpJNLXrTM8ODnSCNYiwfDv7vwOrwshpWh9O6H6uFLuY5JBV2JwwTpUU+94VZ13mY9H
+LZUzFte5yy5cSwJROwchw4bk9ANhpTF5BRXrUV8Hu4rhWgqSJ3iYmuAckvDxdCykY3BVilAG0Uc
nhNQB2XCPEClxnybNqUtI+u6d2vSstQvTC4VPQyCgwHKce82tA0YOkCGPmvfdoVsO2Z8g5H1pMDx
eM7mGU3D8UC3UY8Q0bHwXRgzY/Vhr/By4+trStq3nVbzPHH6SiNxeRH69kpv6OkTotJdlOHhT3uV
MxWNFlVme09t/HECwAydBVgLd2IsqABLVsfOmkWt8Z/A+aWe8PMXQ1FDaAa9x0TXY7s28CPaRszm
sEVtipja8dtJ222PS2gr6UDzXVyBCvVUBPW22UFxwIx9+elwIpagkHKf1aW0szP/w2ieOiB7GDWg
AFvJipmIPvpP4JJTnm/FXEzCWo08yCAx4B3+FIHnVb1iZfhb7jCQT8Y0kdsAJAEqsJo5TRKSmcKE
6ocp4bePdFs1r8pWt0FtlZ7mTgCXQAVle4fx+ESTwO+/pC4Wu5MgT9ablV+rHwPCUuBOec4hCLFM
iCxM0hfBrJ1933mKqf6ycFnRSi0Yoqel2nnyd+4y20PSqL/AQeGvpYzwuS5FbmtsDX59HwNxXI+c
UJMqZGnVu/t+KxUpst7HkBTpl2UP6aQFLt/zDClGYhVFtuRv5wmUXmEiTbxjfpBXyqgEviVwdlbp
xx0HiM5l2a/ENpQDP3A1toq5VGMEYAIvPFbYd3Nbz1n8odaoaJfrZWbn/VKK43MIqsEVGOXpgerJ
4lVswKPgfQ2JoMLXI1A3EMT5/9XCXBOktiR6mGlWBg8O3pczuc6eu336+FiPKj1jCZxGDKVN9llb
dGxd5uNYOZWcWOU7br+3WPW8nBaaMoofUoGAECzMK9s09KY+9Xw1YyAAgIOWO/O0B0oxBCPwnPcf
GgRKll2AJWDnYs5U0BGG8kmhwJKTRMFIUtVtOe5ZcONQviwRRQZEumPaWYwo0BUFJD+iUv2Jxd7J
yhrAWN7wLoaQNBf2Q9ApItxBysp/f1tMamkj32soVBslBhSzJTCFmUOePCuUDEOXgRcVHUC1OImZ
hTH+jQH8uGDgOd4xM4PyO+BFYPHyeM2t9ZGF7AQvnGAppW3rdbcsRa/UHAu3Stukx0io9nnO4QRK
jC8fiZFaFknAlh+vAZkgMqZFoH/w/L0PMjop1kZMMJXOo5+jD0fWu2M24nhqV2hSbDj0aMOytVex
48Mp20j+pn5VzACEpXCk7CmzhoXWZBARqXA9who3sl4EBVszy5uwxYdAb9kyhXfb8byOU1A55suG
q+7jUK9G5Xi7I40h71zuGPV/R3bg0qJHqyCQWPgDg5GRHt2v3xjtdQ8LnnMNANlsYkvpkB4Od4xu
m6Y0ZZ14/WP0rNGGsxDdF2bDsvkOBmQWNIdnVcDN3VDuRtwGjeFPpeBiStAhqPoxV6BNmPKBvUdP
ikO15nn4YEVwg9JGffYpxLEzL6h357tBzj5id+7zdMF6u0vYMWy1Vvlz7n1F8UZ3da7zEZwlD7cN
JUutQtXMkVGGZeVcAmj5GIYkrklBRpGW7oFiTyj6fW9gvOyWds5JV1xuYDRdbursCdgk+W1apcpK
0kQy0GSjtJtnfCm3DB+65DZdufwDQAjHuUgd+jqNadX7yvuxui6JzldRBf7NHNj/dOgpTNiNkJU6
Io/H7J8WdAkTFjsz+wNfikdJimHPNFXWj0VYQ+9JEa7RnUSD0vEHceYb3ov7VUez4awwuJyLHvWt
jID5gcGKw5Gl631xXGBcm4JVXVRTWv0E6JF2l0WNOKi4ruNzrUMvURsnqbkj+26t7/bJOlezN9YJ
iBYvOUbLqwOtE215SgnfJmB9maCyIsRLGCVr0K5u3m8mZEhgvkTwT6GdnTPxghJ/TmSQtD9gpxrn
gL3klTAYimVgwYF0dBGmeswpZtzI773cYqoKFCOpU35Ak5TYXDl0gp9lcEoF8Z4hlNsrCikZYJYt
MmeXC+onnmDSDa/XsdUPRqhUwUO0A1uH4iVvZloSt+yoj8VuKaEjtaDLgz+2Xoo45AdzuGfxn4cS
f2FY4WzZfwQvUGLKR/ZiPSK6TR8bVBfARuJjS6nZ+RjC27kwJwRh7Z5LBZ/aVwh039lcNl8JZZn8
ZPyhEmxMzHjN/JHRenDeA/ZGpHQDXTKBSIOPP5x1dfpa24qwx4kRzZgSt0Lbc9OFySATnnv29xBJ
oIgr2qE6cXvZNaYTrVbST0uanlWBLUY/mlfyi9CM0+PY3c79UECq7ZsGPrKPhGp3PtvaoS8nohLL
VKa7CnoSLQ/ZqDWxINJRrKdrDkoiXRGkNm/vzhNtp6ZFPAXW/XGYn+dprZ1ThLoKHTQTHAYlQJwR
CV7TOPr8/CCQ6jpDO0TmqWq+tYUDUS5JB4F+ZSEwXhoNL0Sy0PflbUmFUdCwSKXgvFaOmaYl8IDp
GoR7Tc4rf4JIQkg+BZo9rNRlV9yZV5spyb1DhQVctiiJg5yNd+35kvUgRHAkd5wEIObMY2746+3U
71alkirYHQkJ5qJOIuBnUlbMBPmodM8Eycnfpb+ucAd8HiEDdVaOoyH2fXHMySnZd/rLGER2ynU9
RH0WB1Z0nEGrVXqvncC59kStpKmuhVv5WQ5+kklBTdyX6+U1Lf9irCTad3tZvyogQCTdoDCRvhMa
bQv6Yyjz90hzJG80WTtv4OnId+AcbQdvPde6TgR/CJf+g92G9zhiFJS3WJykyia449Hw3BPZRWSB
bI3DQIZh4lWjGiXKQ5h/oYujo19PcvT8u6PfkSwMyl1MINT2uoD5yXSL84UXy7IXbOQqPv0PWGsW
2EjMErsRhPxaRFrxT+IK/Vl/eHH6Uod9WcY3NVzJT8AVuDpz/CSm4pSdGWNvvW0T1YXywTFzleoq
8BxJjwSjDPzu6vlvxLgy80fhZ99bbzpP9F6yFPnLzwS2DIujR4MPIVIXXG6HPm2TJ+TBZ7O0thK5
TByFPy8PlcUjNINYFecqIPlPX5eKp2xJUlOnUPbUKlLJzIJUlK659HKFYmdc1PWvExWsdH7A+gGb
7OK225Yy60KuVU1QZrDi2+W3pIC1BpnLaMvMZysoP1vxgaKzJQbPyF4aCld+dxEK7xB9oSAhgh2G
ygtnxr1DM3oAgpJmEhlAmnQUEWUpUfdmq/d2Dy5zmpPalwDrGp6qVtv+39pzvy4pXHJ7M1m/j+ke
08t8D+mYgyGfPRPO9kTeT/YP6cUlBUPsv0mxQ3ecGm9/XFmFCWA9Vf8W6jg9n8zBu2f81rWO5A5l
DGdd9FbxpMjiloDki3RoyEvgUj6ekCVOO+jDUB6QwaHYnVI4mD/5z3H+Xo8QTpt21Be2y0kZXPvx
zKsrAsiGjZpEYPl6CdOZBbRdyAbuSAnNcjV2ZKJARa9kARh+Q3o1N2RI+Wyu7uZ0ZBHsaTvq1Gh4
kWAd58TOW2MqnEtzDRKT/fKBRbhYQE5dbf5Fa4RAlbvTVHPziV56xnX5zMWw5p9CVOCZgnjzKMfK
2MV7BCrC9AU9gBSb/HXAEjtkkRm3NL0q4bW4HIYEcInBG0n/JGAS7p16EoymK8Ero0EFnX4NSNez
AVsk2pHHsjIwTSZnz4ekR44lo7iA5mP8nXTQplLr83E7snPt/i8mPRvVmAGZ4IcG9zZO/1TiZRR+
Hwop2LT0UqQQso+2iVwZ3kfBxHSmRc6tfhhFyuK22myM1viTgRC34WYyiPTSRwbwcuLwzPucyuXf
HfWm0Qz1os3RPVvSpSFOgrxjGKcm0fCdVY35FYwVWq6qmUNf1MS3lgi7fDTmrFmFC9y4lxeH7UZ1
JsDL0wR2ss+ozdP8c7a0Hg7jIon2SZTzgztqHJ/ojd2JTPki+q5JmlBAmlWOFA+IBx+9Qs3Pfiww
u4mhdi7ycICaKJs4VXZRfYqxBcAKwha1eovXKQqHzBgk8kJD4OAAqcGiyGhb6IydO3BQSoUR7EiH
MqclCZcK362TaUWCQ+B07mbXxywvcJnJQgwRklM809mLvkb7bqGFtcNqCUMxss7GdUC7L38oqvv3
2en33W6EqLfNa6LSQHPRFw18fCgpPMpRvq2JdjHlofrHIG9rX4M9cTXXOdj8aN3pNQYcKeP11hLD
89IlEXRkkAfTbiymxr4r1jMqgRS+/phCbhmeqI4lIwnja09rsJMb6ayK+WqTIov0R+qGfwG+vjGT
P+f7Yq80UaNatWkHWl0jblnLB0lbhnKCEJIJDvWuoNT780frgw2R8XHpHLWOTXZ8oOfZQ8m0uwiY
THpxcNhVJ2qX9rAzbaMEHYi1NyzuPQwUAxFKJFzs20VVpBKBSaglT7UgV875rxLRgdOvnoq5HKpI
d5+zgO6cY3uGDWl2YDxphoKiPNqoX3PfHGuOfoQCMcAk8IUqmiyBOo34vnrkRgP0pO/GdmSYCgW7
Yy8F5zDci7IOqsWGoBbdjtILS4hKrdfqaOeuXHD+bpEfWlrhsxqxVYCkynacrX7hth0VF+8dZhzC
zyfl7cSUMbpljWInFzcCnUKlJRPn6p5rJVKtF+82j/ICs805q3SF6MCmpDBci33+k4JWehIpmY/r
BDV3INAD9/h14xkLdvB8KVd6O70YP+UWKmNiBIYklstjY45G+ccX61IsQMGpPNiKsTTfIaOQ3n4C
Khm0Rf0TmSLwq4pqcACvjfsrGNe7N12PRRFsYejFNFySl6CO+BI/I0Sn+fuY2MEK9M0gB1XLcLZ4
quMCnoAGBdjaZ8dN01vqBCTvLRupHnxx7V6s12Cg8dB9YGzRx91bYNwSisWGC6OkbhjtKnQ+yBQY
S4r340OF0aehHr04QPk+z892flHOAdB1DbaeY7KmwaVZpWiYzibmiGfkODCmGVw662wZm7JpE/Gz
fT9ZjNSH28yhqzQuWi9SU9oxUGjF7cdzLFfMHvD9T0lBMbkA8zd/j3sgs0dhAVDg+f4+a31gZJWc
S54fXPFOSDqbxnl4oJEUFNu2KRUiUSZkMuM0j6C1sQB5x4KP2O4t6isNO3BlR04aO4JD3S0zTjv+
m1VEO2qaKpM06XXto8QUskORw8Tvs6Y6eNWSRkMerwahe8eR3UXvDaZjUGv2un+R8UCEwUnqwrTa
EQPfTNkyP0gqK0lCEZxV5Dpjm3xYsCxxsKBstGi2lZrOypH9p1YeK3dqOKhWgp2LM2yYhiNfqFnb
nw7MqRAOhRxcSyF/TD7MBAIdV6hp804/i8v1JC+3ikMtUDwnMhBkq4FS/EN99byVZG3V98aQJx5n
OqYu6dA5ANV+nUxixe1UtYQxW9nQZ3/pWBIEtQs8Z+HbgZkDroV3afdC81ejn0oau3A/7muXSXSq
TPDPtSphIvZF6hZM/8K5YXmletiXUdqyNsr27Es+VzXEwgTv9ofqWK+z2bS9L+Lb6KARSD6Xrptm
yql+pN4hFfhOpkqdr8a9f3Xn/Mpf2v7B9MerKIUxyctL4t6ymDONtMe6EBRv91FneerZLSuDz5pL
2zDA9/K+FLaVllc3evr7RrAO0SrPvWylS5rTjV3KmZoLSO4yBm+y0DtVUmmgDmdBssDQIAcQIR/B
L3rv0n77a7SWvAofDgKL78hVJyIqdS4Ul/lpE2OyOpyI6MHlGdA7lfUEop5gBkWSVORaNS5lldWk
VbtDULX3fekQC+PSW6S9nqzzE+Jbfw28ycGz2IhCnYsF9KiFDSbJLAtmjklOJOnc46+nkAr/F0sM
TcL8XzHy64fcIPxBiVMkasEC5e67rXfmnoVepl0I4M0hRwZoS5Q8tX2GYRxdoBmliK0HL+Bmr8ZT
rgPJl3SPVt21r2FKA77Rd2yRIXV3olC6P2gmGf0sNnCbJKanpy2Qpx9Ck1Q/5HDY/00HJX60uPcU
5PR00Yk5Ipxi9UEtvoywsxtjiZ9dOdnITjcLgAv9GpV3ZBAIU65IdJ4XbfYkP912duHXt2pRu5wW
T5jgc3s8xe7Vsu5mnAoS1Zb/T4RSPOWV6HI3Ko/kskZrFRutxVVl1GIrC8HxmCXdC0ane8iDajBD
JE0eX2NaMHMQWcZHQFZAl1ewLuxuIJ0qcICaSvuE+FVGpNmAN5G4i1Suy/Db3MuCb/B6nogCWfAk
AclYKvS6lNUYZBGAhMxJFKfMdUn9jIQ2WkBG8icl+nU+1W3gFh3fQrPZwhBAcvAMfb1FL1kiXUjo
EMFtbMZrVdfeyLM5zwEt+JJ+MFDnhre+eGqJg6b6+vS9bSb3LmzAokC6Rv0H44SRQ4HW2pHWLQl6
eaLW0Mt/1fFBXnBL4bgv1j1E5SS9rxugOfPlwhoum/v8GND//WdO+LLM0sOS6ereSo+/kKdw6Ip+
5kknSIZgpMeK/p8teGgUHfxIWE9sZbARFQ/igkyB6qehLU7sRHw3G0xzcXUBmNrfRm/jWhYjpaED
ilL3wp3IzJHJUE15VkliXFQU9XkyYQiNB1IbA3s11VLVNT3cqKWdsQYKZiNRImUHzcmJ7WvHRM56
31/qKMw+8HhpvgF75YEFHlhR6fpuc6lvXh5ncO833s0p4Wmx1VnYm7fWx3e0M71h3NtVoMwVa0Ge
DOG7laX46mUe88/62K0r1JtAxDaDsJIaxaHyU4lpsr4nDg79yGSLr0YqkZDuAkvyuTxZ+IgD2/YX
D2zdum0hzFmqkobHFVpNb3/hRRnW/OFglKLHyuRppwSVYXwS/VqmIPstH0idkyqoW/kzsGggrkn9
hCRVoQbWB0xuZPsn2X5X0BN4KOXIxHaszQa0y9p5LyUUrGZq0We62DueWgAnx4jR/qtNEy41t0/I
PQy30CwBg1vFDBLkusH8tQbih7IaUPrzSNPimZOTMZwYOuMgpJt6Jvs4cOQV9AYyDDHpjyHBfL87
s74bBuBwNLQoQBh8xMIHwtzmFZuj7nhSUtqPXd2xIeYdWO32Qin4I8DBQ0sQTfOqB9YYUb+CV9AO
IrlJX1COfbKpyCzd6ItBrZa1NXMaAT+aMoUkesVfxS136Y614wVtYnna9imFe6x6ASs4iIsnNalg
2/XtcRUh+pOK2YEAo1gsQEwV0pRl9vUQLJtMNGrP6CSCFCq15GN3wdYfIsvWIuUBO7PnezjSwSbQ
WpSO2U8prUNpICS2Pfi0t9k1ifp1ai+neXMJvkSKzsXLTocjewP2U/itLg/9qcxEAvq22/JQDxQd
YIDFBoHtUTnfFiU5gJDek3vUUZaKii/UEdRC7h7xYh2frMGgn6LS6C0Cl92T42/GG3tbwZ3DVA64
2/IzChO5Y4luFtw/h/IZ157+cOh3j0rRr+NJcNH6KoI5D9kMCOsw9QSQhaGGhVDK+UNEDu1MRJsA
XTxAbqdDY+TnKkVVJKU7fUg6TD0DZVQifrxzfqE0Y9X5mOxjpL54GEYZNkbaFFXlFrPs9RAK9AZa
jmmglIiLu3WbYkVPiiiZ7B9DfyVSuQoFl5q/DFnstYcVb9vEazckB0cqxeS2YTbkmRe2lUUQC2jU
rEA15uDtG5Bou844ChzAsmr1z4bX2PA+RisyexbKcrvobDJBNZogUU0YSOtSe+D6CJU9qb4CThVS
T7krQz3ssqiYuRWXDGoVR/IBwFJodRWV+DQH/fHBUilm8r1fCDScy3NR+cqUvbefDG5YedlkXEkZ
9InwU9T+YwFieQJU3ufW5cv0/qiWRfiCt+SvKCKIMXUTCjfvw4a0mBpHSHpybVjVDAww1HUmUvcB
eBRkgxQrT5pnzKrhnVWwnSG3DH+7pIbNKIp5oJ3l9zmVhuykf11slw3GGXAxthRuStHem9X9FjX0
VW9vLzONWK9JJgeExgm4Q8GZbmYw19nLj0X+m03cnf5LFqfpL2dRydD8RR5wYCkry4lC/hFjGHIA
CgXDBabtmKJqfulg65NqE6rd45v7IalJWXYQSbCWotvuGeP4fTdWawM25mNamvuVj/EtaygrJD5e
dyU1p/RpgZPfDnPn1jjuj2luKw39kKLqBp1VehEKz1wm+V5V6oCc+ioRqCLFNPdyO+q/5YO/OAad
LApqRZL+UmMYC9lFeaQZWSLBlXGQut7d6Ld3TksV0bAWOouSfgGP6XtcJ8VzV4tz/W7RF4Lax1fR
QmCSJuoOPx0hVAgU5af6X9zS+GwvvR0pSaxcem0EpdxdDWVTM4Zq447voIDm6FaXz8cnMx7aH0hA
a06dIgyUExKg927reguNUcQuyP9qDYMG8hzVT+O4DCjMHxiSCOsdufFyXMpq/ZwmF6gweK0t2wU3
mjlbSS13a6MHxEDpBN/NUSmGdeFQILCLFqyvrK2fBN6r2nH/YmB3nVs99M0Gui88i7slVrKKvgVj
c1qJGs1sMaFR/AFuUIEx5guAvj3T3igOF77UTYhpo+Oc4owqwM9p2g+6tgevHsEU7CKQURQWmDMB
h9wsmxjL+SOUJSy6h2NM5NZoHJbWQa0r4M7z7z8HCORzCT+4GyW/Cnad7988TkC3u/tlEl9DbrF+
Ql1WH/hLJ7NCt6bw48+nP0Hc+WaWVhDRBW8QiID1uQrWvHyV2cbjqcbPo68qK0gtua9oqIR+zJrx
t4lCStAMBB17pa9fGuAW80Pu/JjzJd2EI0u3XulVsnj4RLvubbRLNVij0dFApSLB0vbP5NxYiI7K
o0ute3C/26vBgzXJPEoo+3TBCexdD3U6LRGNbx47SVrbJLX9PDLQF1s1anyCkfIxDJDT3qaJrECl
4eGrfBigVUWUhDpxQme5jajGlpwUX+rcYqImN17DEBOGVSIu2r4eo8QYeojMxUImauBdejXxKUIY
n2VhZ0ztPk+GEXLrb6NcI4SjjUaqTxSyEl7fg4f02U01ctIreVRDynMtJ8EBH78rTZeYFRjB0tD1
rCZReDYqa7JgnR+c88qwUrNDU9LLUBdSJt24pgBHkWAqOMLQeqjlpWPK3q32qJM/lgdsvcqd2eg6
6aCY8fcWwKuw2QMs1TLg7yVUzu4s6e3PWfGn3Whg/g6kQhl/Jy8ny52OmXBHRzpqsCPaaBmYSa6F
3ojYiPyFrtJE9bD1qNtGkzTKR+yqj6t56QtpTcJuTqKCf1GT23NRAW/RdT5xdf7xmyZV86h0i//p
bDLPweMsLaBA4U2GRKjMtXbplyE697/I4n6A2Y/74kNI7SEdTnivYvpY/NvPentX6p1lY5EBp3uD
QmL37IG3Eoq9kGhrCCZnOHMRZjWWFljN8ZRzCiCQr2Zux7XBSMAQXXiSl6DojXUIAAfGiIfGTXuX
H9wYrjX8VQ8A3iaTNHwk3MpEnauxmfbEZYC0drDU6MI1fx0NtaSi/KPpCR6LZ29ZZMoCbVoQewau
QEftN5fRX0iwbt9FTgNaZnLPq+r9qqIlXdlplGQ03WUyKEcNVTBwMNsLrPzq5OUayd7q06aX2En8
DS0iEt/YLSimD451y8yM0peT9kfsTdJ9QvGiSInNU+T/0+KtSqBVOi9sPOMf274TlMidsoDTF9ML
ZOgiPS4czkEqdQtvqD7yMXUGpJ22WORpDa9FwiXGXPujFS8i78fK2nwtf67AtuQpN8aHMZ1ROeGD
AI+Iw2YCmT7W5Wp0HECdflwqnbPc6PPVxz7az08ajbBvVVMGUytIMTrIlTVeANO/42pxkkNuCtcr
nA4c8XcT5qmtoQqM9fB2eQpFH0ZMbUxL9BzFBMyLJlazUDrq01zCYoOv5GaBwvg6een6CRDHZXM6
ZGeVT5pUUYQEmDVq5pGqxHwzEzJumz3PX/wOZl2LUT6D5tP5a0ZYQZrIs8coMM2CjF/dxmPtjj9R
P6l3PUZGwG7AIxqfTPmht2wB0rP9qo1K3eNes4R2/XE7E9KXETL0pG6KOPULrSbzHhr33ZeY8Ye6
KZJc2OW2O5a2Vipm7YOHPx73X4dZNpf88iaNSRmvLIKYsXOzVWS5h0nSgN96peKlf3rcPuPMMxsi
K+N2n5TH3uyiWHXO1hplSf8ZcAMSMVcT2Len7whpY1NG3jClUGH+gJlwoI8MYywhSAHigUFi9myE
yBMdz7K7tOSB7OXFEmkOvbeuTH16sQaJ+lIu8Nmez9rkhcDlkPeU/Xc3uG3hNh6PXxUqKuHidwaT
pxU/WM4ak0pPkAVd/kdjhO1THaXZ85WxgiMhRu0ON/5+bg2CHTBDv2BaDgDhQHDIclIvv5Rxtryo
xCg41hBwdNoKtI9kPahouaLm9wERKjWt/D3MyxtTHySTNWMNVrEkPvb7xb0/STWRJHJGOGDgoKC8
BCQ2OShcPF2Zj6MRTTlD8mYPvx/R3WTqW/2sVvN7VsDf8IbhX9Tbl1DeSPlkpGDoUyYsVkBZ3CnT
0UeWdKoMgbK11Ct1nbc+JrYTjP1+QiMkM2bhU8GrrU56jhSwRDxKpkAgSkW/476vLJWnGY/rqhGl
Zgph2qEzmYbzLEOjpT2oL0pSzTRUXlC3bYHC8Tyy+Qmyow8aNVRTM9SVCO7CtBy5j+3xNy4YZXuX
e5i2N6MCGeq7RXHWr+aXWuCiPcY/Jk1p8k8NmU8jypDM44vFP+bXHcM2D0GmSUH6AWjdB8zue6bV
ddXsxYdf+3WJ6Qk4+62jgHNLxMaMKDKG049FIAE52EML8d6Y8Tf1BjVpXKZ+HEU1iUMUSqJNVrz9
QwS3qIJ2LQURH4hJnva0AKohBVi0HxIW8kIv5HwPa6kN2qt79lEWUKARGDICP6bdtMY6QkraGDOy
NIUtw7neUjiEp3RpxhePgGnMwaRmtJPKMDv3JZ3Ui+zbvV/ZUfuxJeILmVjRGAg0CVpfzNRrFapj
RTGQttLQ25Bb7wHopX00YHRsWaK4z0fGDtwQuakFEYYqkF25B1js2876Vu1npdnvR7+YTsdSA9L3
46/r53IgqqpCpAT+p6k7lpRaCunDohVo2BgNKKzzDoFGTWjWRn303vZUBRmwuqtVFSgLZIM/TGr+
G2ORu/CxjeNJU3vxvhv+EZwWehZUoYYYO5SjNRz1HhTCuqOj764yNE2UMy6DXon6ndh/mjhT1y8e
7YcS0/otRn9ZVoqAB/KTpjCOs6W9z4x2lTB3g9MOMtHbNXhO4nSmfA6wmtWkAhMqab9bz9UpJT/s
lvLcHA+1ZRIMtKAtlLTsUFi+4wqjeZ2R0aYfzaTZFdt99RiZNZ3UkEXMWAGZnoyAKmjnreOK1JHJ
bfrWIFMPZXjOZ04BZcbxX+cJ1jsoDwYEqRkyloR4U0JktUwsvCBXe4WUhrRFEYUJaHP9Jo4T+SvA
PmlCAjd88BRes10X8S9faj0Oju0tYfZwLRrluw+msUn5Ni1iEONouqxcHefvzxW7Y50jQ14Wfwoy
yI6PxojoT+a37yyDhr1+pPiZ3jem0t2c+32q8/Nt9muiPSpZwM3y6ty2NdEnfS/FmNw66lLtD3u2
DVjVkSbHY4D38fcYfi5He1NZ2p1vqurdwS1rHyoMsz826XBsBuCV/xu/YhN7vuUyUneTNB34dVxJ
lcCA9TC0MAybe/jFMtqRWL0TOKkfaTkRQdxhmGuVi2RQ4TZqF2JyUOSmAPc3l5uSyxlnMSfSPPdK
YSskkn5YeeAy3Jo0nWkIiPP40QD+8vIF6WhYPIOH/6zgivEn3EJvF0ACoBUI5HXxde3oYiJT925u
pumLtkJTDbHmbhmHuJnkLDbdz39TOFlBICDNOzr2urbvogX69TmNoj1GGj1q237eh2QA6NBo31um
sHZrr38VqlEOgRBJQtm52QXkesnit+IdDCO1M0uIhXXAmTkMJHcJ99wvjFBphngqb45t3S/axPsi
wJk55jGLGn0VhcCorYQ9LbS0BILtViLhSZysTk/skU8cpcf01vRB1YSuzS/aRUgqBTUpyeJTr1wE
ddjcrqIK7dfT7NkSKkRTFcUt5ZbEce0QFj42fPZ2FCd/z6ia1BcGR+7DOUxf/iE8ZyqEF9CaJ8Yz
cnC0piNpQ8PRVbUgX1TCyaPW8taSvdLEfrD1Y5S5XPe5J7rPNzgSw4QVCbd4j9P0c3l6Lr0mS7KQ
REl2G/btRsg97DY1JMP20YDWC4hA28nyNJ9gzcuioDp/N7siqT4RqlRQ6TqNAyEVEbpTnSiC1oM6
Pnvp/uHiQi7Tj0mMGpsTDKLmhdq0aFu+QkfezGldRruhWA2SurKGSC2bwaRc0BtyfuTj1HrlVUmN
lBrzHEcXFXEliBtUad2hqM/z5EjG4mfpMycCu0EQYM21imSo76wJNIvrZIbEXdTL5tjDXtpng3dP
t5CaRAHAvrwBXv5eqBslC0d1/M8pHvQKRRs5jOIdn4Q/vP0hp0++2EoufAh0OwIT21A0FMHSzaZn
t2nya3GxEJ4k6R+InFXSwZKEhbrN83OwtPpmFNymTM5V/1oHT8YNBeOmDOdAiYePtigAjNFl2/Zo
GsklT64ZAiX7LcsJ53qDpFn1CNEkvX6UEWdY9RKp5jZ25ESkKVPmjo8osEyC67e82aOrMjo30NXZ
xQBW+0qgrLuJa4WLjl10Dp+omY69RpoES9bB1LwUnXgB1iLsTtUq3ken0B3FjDfsDIOjz9hWeEsW
urrDPqt3blvYMezaA0/XR65QNSgc4+jH4yL3FKZWAykJRX0/wd2D1fdr9q2surcqPJ65iUzVDvpT
BYL2y+I0W4gF6YBV5LkYojEyZgep3VBtDJdH6B9mhfGUWpdDy4ppCWPDGHxDMi4wInKVRqJgYXje
w9kYJG4P4UNpkct741baWKHIFox5tawnluR5hE9v4jKPuS0B1390qMYDsHRwEJA3TdmrGM5zkIMc
Y3/BS7EFnp7JhrnIY6IiOIrchBQJ/V3iTtoTJ2rVR3onLBp2o3jh+2L2ZECg7VGBSHUksSM6GLEJ
UnzPdcEJ9kbi9vNTfxVLQCqOoqvhr71QdN5y3f06gVoJ6wA6LC7YOwQv/ykB4jQLOxmduNAs3yt3
MvlRKDYI9tgeiBu31I7EzCv2laiNlHDckCLgpaZiaFE2Mmrx6GdrofoHnwJevPfcOd16lyZULOHZ
zKhAhzvsuQzNCAv13iq5cBCZVHf/xj4ly/FOtCLAkwnvHtOjJUp10S5tsuOLWrmI4FG4LDSrP+J9
Z64wveNpozwk5xKL4Q4Ad+vxsWcNawzWih6QcywKvigz/R4FAxQ1wN8oJsK/U6xeZsWXtaNmSNja
4zis5Pc25x5zuaqpkFCHMCpgWPdxk7Xsmu29ferZD6adXCvhwPdlIBYYzCpx8YalrOUSnjiXGsXb
R78KE6nng6yBzy5Ow/iytPt+3nwthewVdgOpRf0U+1N3WHa6kdyiG/4p54elh2gnQsEpHoJkhCDQ
SDgzm7R+AQV5BJaCwyariBNNnIxRpntn4YpOctDaQjjOb6oT8fME0l8AWJIn73QLBOMeOGxYeYO7
aVtxeTP2ObOefZaVcqDK0mJoV8Mk5QJqbQCtAFVo5v+dXo5ZNk0VoKFGZEGtv5htd2PKnFQAgfr1
WInFn5z7PlrgE4I3EuAUL4Qh8JALqQgamiBzwDwtwGtouMSu15GtqMSZlZDwpUXLHCZc/sd3D/EN
Ee+fOZweXB6W1HPcZLilxJcL0Hjv/tWD9cbzGKNsXwliOvT7Sa6J6mKjZw9YpvMK3oRBj8r0HXKX
z7cnfbi0czBjJYh/fWlivGqiXJIqRt5o0BffIw98xiLEaQTroXdtLvvWKy7YMmCOT9mQyaYlGY0R
5QucrZDBYWkh1MbtafB1vrhzb4ZPiyAWYCBzkzKeLerTu8v901QmhJs48Y+ZaoCkIypY+XdYWaQe
swyX6/qv62HB99S+gfrYytGuOWVIoFm8FCzH08S8YVlrdo0Y5+aACE/JGi9ZHAJ+MNelP4ZttgIN
x1gtcNqsVR/PRqS35Z5YYd3EfNXXsdTdsJp8kWQsfECWk7TORBKepro92rM0qggtM70r1Ndnh98O
bsU4nYINtu5AebKjxwUUjbHmpo5xxpRP1XB4u62VOf2NQfVv77NwhIexXs/mi6eM6LzxEx1Zeeui
Jd5HsYBrzqrxDNRT28aBjqxVszCWGGcjg0oDERqGbmrxHnaY0lroG9ugxwd3MT70Rds+ZOw8JC1T
gNZxlcjuhTd0K3zTq5ut8B3uRWwqJ/44q8jc9XsGUY/fUQ63FtSU7XBQg9/5xvUZ8giDoq4oAv3/
cVXC1U6H2K4+CrrXvMkKm370vauHfNraQa+Qj042wGLZ1x7qQlCViQAFNLQ7EN/BpBrd/7qvazj+
aVPzsX+ftDtA3YOkPlUdpN5BHCBAV2n0GAn+xK7RjjjIruGI36P6oVHLr05uNzL1neo0GwJrnAID
R1yBisO2wdnCmpk3QfzSPW8vsTie8hixx3UEZhBDIGVJGOtBR6FcW1LoAIB/dM84ZxwB9zx1lBva
nzanvZs4RUNbLbOKLEkaFAw+sDJ8alz+hW8VnWds3wnKI2lm2wDxD/rGLvCSJ2e7QUZCuIIENiZ+
dAESAQ1C6yWo5h4xWvG62SuojTmfqHyGH/+tlvfbjbLM6jxvssCwNJospWTJ5JfpxE3NQm75Nedm
hBoR0xvFXlEBPdJkQboHSnOOvZ3u5AoUr7iewEL7XB8KRAlbc/p+ylittHdO4La0YgZeKpajNUVF
reRcL40rxRVfdRICuge+9o1eKiSHgStW3y5uaIhaV99Z1CL2MsqDXi43o2UIZUinyocgwfrwI50r
aegK0zcFTbhuaj/yiOzZvvcYBD486NkCafvyU8FgB0R9REBrYmcIk59FWb7MaDYr4+7mpSU6Dthm
FNr5p2sOuv7zn69+Ta67kGoIWcO9FdSHkBFVCweLw+Any87dZbU2VDTQkx76krIL4gAbma1/SMBe
wfvlUrOYwSPcOiNrSikAg9cJi4EN6leYNTKXBm+664y6dxb9itDA3ixfHGByYpcNu48OZj1VVvG/
/2zA0gBQ+7hIW1Mkzo8ilmpufvEKol3rzqJFBVYf7S6AnHx0HbvqQfsdclO0RVBWP7zhugSDeUY0
uiH2L5F9FIoGuEG+M/Q16NzjCix7pK8BcGRujDCGTYacL21vbfbibCoGwrSkJdhy9JCwohAGlD4R
KpXNxwswFoxMcXGv2YUxJ1G4ZVuQ17aPheN7UDkF9v5qwuHFv8KAS6SfEUOjtmzOMzLlGv1QoDJs
yfbdvxn19jWovYJwH/G/oEeVJrnXo9PaCBlkCnIn7tBwKNauflTLXbnkE9ue038c4FOdqebjlgNd
CjTLGzJa1nll174/yRVB7JCgqDnT4IQXaT3U4r4TwBxZekMbbN8NIAdZ8j2coyEgwdmTF8pbnNM7
vZgw/v4FVopkXOR0y57TE3mERDEG86TPNM25hfP8yo9aFhKNykZEt6hxLv/JItxYo0+rrio6SM00
yLy9VurC9d/L/xL6kVG0V9llN1+l3OtH8AYip89cxHqVmJvhW9JSYpg45QXhnupsLlc4oyC/5/i9
ST1glUT9vbHfyqgx+aRz5VY2qW33bElIe+bKJHv7UmobvtZdn50FLY6wAKk/xmjJ2/wkGPwYVl6L
4w7bSQIWGT2K4NPsSB6ypwK3qF1/5v/qWvJJkEHiuyq4GS3/yIZVwkertMFKD8XHMF/smQ3TFKxb
qT+IXxQ1vlOjTzW7Cnp0+MI7cBmJAxLheqIYtpbHHqV4qgGs5HgiZEQ1ZxRZ6QBPYfPx0zF6Nbve
Zp+RL+2kicyAM6KC1S63ss/ZdZxGk3t+QZ9K/OHJ51Jd/TYRqbueXJQ42tOLTvuQUAkBGg0qa5ge
AFTPOV3yC/ThFAS7DjVnMrAsuwP6CI2VgR5ChpQeZx57Ou/Suv97ySzqde9z08MTTFCr3FOonLMD
C5JIDgo1nd1LD5bDmEAClu5tsr9Q3UWpxdRvnI35oNuNXLrOlhuukThxEwT37tldBxhpPO39oHGg
vrQS6KtEqFQ20DJoBRTRLd8VxLx/fsCksKlIc7Rso/k6gHm8lDrfAbp99p4bxU/vt51bHXLK9beS
vkQRvciAeCv/omOBuKBXTxzsvFsT89QxeKbB7JVbUUJwA4MjcZdH1s6dDlo+8S3xXsit8XObt4eA
MeH51jGAWYSVh7zdFc4RYVW3kYz7k0DEZhaVVZW8NP42jlFLbaA3AUHI1zLJ+ezhhv/tbGOFmdXN
u15Jp9bcpx45HXwqwZdEsNGTxoMZz+65c7NPldUwgeuHiGxLjFU0ZHSTsG/F1H53HQgp/zZXp5bf
N2GNruh4zhQ3BPDPH/iQqwa4GaPnMGS8yeHgQOTlAirshYoEeYMecABkUYyRplJXC7JQ4SypKsUx
Q+6awe3A9Dp9SeriNOzjaojXhPVKq/EPDJck3dFjj+FfH8WKEDYllDzSeIiGlRuJx1NzVxhFvLwm
yCIjmMOKCTc7RYCrT/ro9InJbzFZuyDCtlno4LVGwVtq0C6N33mqnwDMdcXIZHBYgSWuWf2R2kYG
jbnT9CNrp2n0hIzmyNJm9dswF/KDR3gEysulprivGSvPytK/xBJ/wgcv4wKvEP2YojWrlyeo6RC6
DrxiN1tWru2AxxT1P0ggpiVgloJ9WMWSmgQpKfh93vYlOnOlM1e/dxDC/OkyK9NS/0zfvOGB9dCg
h6PgG4dn4aOILR6RCVT8nHA63ntipVVg1JUyR+gLpBz6h2lf2nXv8AaGxvLbMtPKE4D/lWdRuVUJ
8hPMo4L2l9Rw6bYmVc9kLbmzd4wy6QWQ6avQ+D3FoNvIySp+mmCyelxCmYdBBnUr/E85Wf/VjBZY
kzzJecVa8Xbn84YfqIWguz06u998/vx73hrHDhmteNHll8vOD4MI25CDdqkCV71F6TD1Xf6wgDuH
dWkcL/t7cfxrm0bDu9ZtQpF+BwarJzclb8IaWp4wxh4PKlN6QLfAd3ogJp3UB/64HuJguPBFSZz2
OTwRtm695OKSGx0aDGIxrEGV+TGFziYBMXJk+nGc8gg2yuakbI0sDYTojtSqg/uIEW8Of4C3XgMp
dNBdIvxnBNMMn9eVp1jqSUzl2q8gIOk0osWh88hoZRjTDgTryqRffQ9EJjKW3DEKErVVaJb8+AIl
Wqa96MUhyV5gm3w6Mqpm6z0pfQaxE1nlf6SardBR9ei93ruCOJfWXAIEarcVXRu49Y0ojlZk+Onb
FIwZuNiEUrZsgeUOuVdRCBvy1ZtRyZPiuIU+prJf6J525VBRxreaYkU47xi9P8MVBnpXwC21G2Di
w7/VugYnCWxoLlQPEsbf+Dt8ze1CyYtjpqdz+4QejPzvycn7tmrnv+R0ce/lID3CjPpsgbImfWxi
7T/h6OHK6H8hTWlxrZJXMl7lNCDAKl9xQzaNYZeEbZ7//iuSak104KKh1N0Mr5q0jnyw9kfOjOTj
BLUuPXlpZ6DTQHIhfxOvTxmm5u/jRmWkvnw6QjSBb1tasHx4pwAr8Yybh3igrE4HWlUK5eS2umcm
ki4F+Ee1iMadMEJProej/CEBNWNFK2us6KxQFMkIYRtATNQW8BpwNhhbVQVxRJI0+kzAbnMAHofO
eWIMtTE/r+sB1sCKBT0firjcTXg6gqWabwZRuysit0j1iNNrvkbOa4jlu9bOB+RRnCE3XNaHy5MF
sNyVvxIqXHQYVXP1p1F+XI82ED+TLx7yFnvjfDEnDnSHgZA8DntmaWqncJ3a8bCCuu7N1vuNevsE
eWbz6Lk0zIDcRWmyrieS5Ydh1YSnMuk9S8nzt22975T4J5hRspdXAriCdA3VC149Ro/G7rHMYJjj
E/uFO9w2sK2//J9FBaf1fwq0fAEOef1lQgpytBPgFO6Xaem25QuI/cfp4O3NDqYbyFw8TfW+DQzF
m7709u9QXQB1mXEQOUW+XfVqBstL3KYRPxXb05RkmBCOF1AFguvAE2fJHK05nkNYrRnPAs/w+shi
OuqXbxCaSD7c6g5kLrs4NZhO64bI0xGal0lLeak/hx2G1kdpn3kW5pOyLmv0QJ0xvJIyrMZLllzy
IJyWjeeRVC2JbHfiW1Hw62nPsxzlNYjc/4OhXZNcgYr+uJE1DoGTZ7+DKsMjc+NSpSAZm6GtcBtk
vs7cdITeRMa9WvEos8ZrMCpyw66Xy77z+71N55L5JKoXQGl0lzPno6HvnIDWyq3d3ZuQXJZ/RoRM
TD2Eg6apuusihVUcXZz3X8/zUKS7drDvkHjV7gP2ZDUgT+o5OsLKCaLt88ID8OOyfFTzJppwfynA
mnjCZL7MiLKuj5YIpY1uB6yAADW/Q3prpb/ZxnPxYSnHV6xcy0JJCpKz6ulL9jciUvcaTguMp6mh
8zq2XCWOOmFh7u6SsjeEdt+8h3vYWwTKuBVXULoLlmeon+2WBXVHAkirfAGgK02L/0Ja3zlPdXir
RhcxlU6/KgFrg/CDlYTJgNBNTqDR6cRr8SpbyZiDmZuNDG5cxkqvOqA/HEwmspeoW6t4IEK9IgRo
WBjw6uo30Fl2laj3uEdd2cloSFNYweZtMpOUnPJHMfW/Pbwkl+ocbcrFRLM8UtROhXM914852Kwx
lRemAv6miJbli07HFvjSDWZosIK/nzghhxDdXkMta6ES59xwSAh8NAVzKnWu+MEvEJW3JlwM9qok
iUJ0kume92aqWv6C3M9dulyB5OhqjQp60Tucu2dyBXP4MoBgBx71iaJvsWuVteClmwn6itmOulgm
SBmC/2OaMeKvJyGWYCtfaMXcHCX5NRb3R+A/kRQM08tiCVGTHre7mCiSJNCXwXPJgGRE+yCotWfz
T0Ah4OKfMYWlofz5pKmyxgPw5KZWu4lgo1fa1V77mxx3fHp7cajz2H4LlhVnO7/DrlEH0gbhoO3Q
dcuyjMuo5iji96gDqY968waJR1tGBy8ia6sB+sWGOu/JAZJQP9FwQT1gM6fzEfoCqcDzLEoQ70gu
01Wi9kGyHOQTeB99zs/lFRy3Ha44kvnCVyZ12vH9n/0Gw2VNhgIT+PzFRQYWJTEXkwCOhKu62fDR
MGrHo6ZF7VOvQliehpkPAFoig5nMfjqpErZtui5ht/7U5rw/UiDYjGP749NvPXbiaSJHs6QbV1nu
6FS717hk1pIoq6Fs6Y/OSRgQwYqOa/onsaCj+xgRE6RCkkBmrtRa+4NdswUGm6x0bZvFwIQ8gdCN
dRG/cZrCNVvrR6ssbDdvUKbaZnLie/ow9oql8YVTtA670GtCX0E9Tv9tYDSwvrYCkawxADtr1E7+
jv1tNzAPpB2Nv6g0oSdIrzO5NWzns8lc6i5Ng9bWoiARe+JQOy004XbnNNB28XomtgMo/c7C3x0c
qgi7i5efrGhfkaGNDddSU+PureuCh+ARHmTjP3BFxGGRj5AdDyIp9t/tecUPkGdZBF3O/irAQDtn
QDQE9gPt8GOdZ2YPkCdDIFPw491N89+RAnmsl0ewib4fNWhyD9jtBzYYXFor+7S8jVJbeunX6GbH
cI1N5EFGFEHBZbKRrTFDfGeZ2jvocQ/qz1+XYG4ig2nnMm6k3M908eSIQqXLa2hf6hbjt1F0ICKT
NwhgMHEkVYGU5atv8hZlfjFaZHIt8m+pY2p3cvFmrIRgJ+O0l4n2FAiL/7a0tdF+Yl6rtWladaVe
clNBIqddc6NC49jho/st557USzJw9/C6Uu41WbYZGPh/W/lXHSuppoydTdkR1MbCDNTmRKhM2ywQ
AnRiXeSbJKwNYzpOBM4tEy+9G4lsemuCIwvp2H7S0qMgz48xAOUQRFRMYRUZNIwTWiHS8tmw+6Gn
1quJ3tKzavuOCwNbUdJ4C7Itl8d/SmG1v88/WGlY3ySPmbS0adxN2ut5etE6QujeEyh0c7qZNoRv
mxvnQ3AMZI53A1dkQkEiLPTXf5uIY7A5HbbxmG7R+EAMyyjK2yGeD8Dx8hEUVNkbuSZFN7WrP97S
bbaLAQj383DCsuyTTdL4d+ftZpi/JjAegrVTxC0V/PRJ0rHAoJw8X6GJik7PSHmi2pmKMb5GznQX
o2pLbluCcRPrDHJo17TIDKcp7HnnH8tV0CjLim1P/yHNTG68GG1xtv7H2fqDNPxAq5hvBu1ePrcF
z5B+oCrRbpkMwG3+bn/XFW5yRTeCosF832DkECHMZGJsKO7OYSwKUHiv83+TdV5qRsIvBUvdq3zp
B4LXuAdyq7VP/hESN2KKOHGKbX0b0Eb144M0YdMAsIevnEPZy9fiGVxuHo1S/FPDNc+NZKflIRLA
axbABL359WYHF8EW7KENMif8sUutAkfbgdh6g+ZRil7pijcP6OvgNWbkvIsJtHUEUPwv0BqgBU2a
iliqMYK2p0dWtJCzzkamrnZ5er1vW8rDPEhB0lWMUNxaN0Fnm5DEdFO1zq8RrEhg+nYaBeKWoyRJ
OCAQ8K2GnQBFsiX2zTJk2AHw2sdTEonpolq8DP6gJlxvjcoUB9i9+6DeLfPfm1FpEUNEyco8Af6B
BInjCd9o3s3eR4eAX7pHLjiawLc6kzUnPkz8Ht4LxcFJenCTvkp7IamJK37ulAAImIKQ6r1MgkdQ
N5CvYfg4nNwpPk/PCgb81hphM66RTaOwVQfnpuc+Z65NBhmTKZ1TRfbV94+3ynTkBpACXBcEhzvW
E0Xarr5BAqTDe6mR4x4ePyJc8Nyo0mbHVeuR9KnXjZl8SfXxNn0xMdoUbgTcYvlMF970x6sIrTNK
jgMjHZ7lqmWSmU8EU+ThiqLmnA6R0xotj5kYmgxi0hpk9HjDkz+VJgdNHCViWfxxBDTvVwI+dXJe
HnqDXLq3TDUlUUusMWKHtUPn0NhVa0nGVXDnZvvJJr+y23Dr655gyCPlm9o6L2ncB08avySF/4Zf
QimKvwzT8S5Lkg9q/4XI/wbHF15eM42X1CdQIpdEKPdTWrMLvQIhjVVpSmdcmjPBeY2XZ3gABhXj
PnAnLTptGaA3lRyoRPTy69pKK0KBpT13+D0+0OX0SKVdIAHLDyOVq8xtZdSDvjA2xsGpNk23Z3ip
6cT6+nUTUN4gqYGqoZURkLzpaIP4dNwcf7xbSuxiF93Te1FdnKx04rv+bInoPzijCO0zKCJa8LVP
xcyEudIuzMeJE+4v7FN3gsF22lGNyM5U5aHktaEQnW5v5K8txbHukvhdPx7n8t23uFF/bhuc4ZnJ
DduooB9a40Ky8Jqj7lc1RcRSy9dRnEu9kvTx80Q9F5v2okbMYoQLW+b8IfKqZLty/AcoNVoSVQkp
0doTc2AgiXGJJet8IxGbsDOTGmuAevsiE+0TBwanVZrljdDBKO1ggahi49915VbXxZApF7afdXkr
Amrb4t/DiSZ1ExmgYbYhZo+Tp4i/WSc4HiWv0Q8stm1ZV/i0M6CK3X/Lq4k9vc7vJ9d4tJPGdowD
+F9UovZjEBW1C/NwrQqkGsNZno9KTPxXj2WyQwDKfq27lhbfMqZxEpt04fmJq1uFJ0Ex3g62zdS3
TwZgry3E11KFM5e9KYIBUdxQhfVcJR9FO3mfdQBWjZfPwdID4Q+GiCEN3FAVfvZ1W9IoBHtmHq1F
IkEQtXGyLerIoH67xZmayWH4Vxv0BEpN/m49/B2eep0/EqTq7v5XBGX7Tk0TkDSp2DY54/Z1dN+4
Np9UFLUVw/SXHvmv/QWjp8r26H0qD4UEry1LCifzGUav84IhOkqPxmNJ05WkHOOWmn6GqXyK1ZEc
xNfcg+kvwngQ+zNLu+BFVzyxwTGNoCV0SLFYXhybfPbOdFWIrlNccLMV24Yueyh0ZKNCqrBHCQ+w
xLL83TgKB0cEoEmbt+0QS8zOmMJt1Nb5ub4sH/Vj8HlcQ77CU7nFJ2UqhUfZ27hj01KXesgIdOsC
PwiNEomk3hMaE5J+ptySwaTBg8MhWvdbsQL+l5+sru04RfFPgjZoZdhxGtLcNKYsIuRCh397IMpD
Ool90NFsoukKUevpPUAsCFfCjCmCtQdrhMBf2KcCf3N1Ub8Fh1ySKlbxwiOb1QyNHbV6/UAYki3x
ZLr8gemhxqtaR1WTI7H+kPl1bcE4pMURB08fYmoQFtjMcw4RcBG0aEUw6RvRIfrQKQdXrC/T3BW+
ip447+WcdvSIqsZQgPibCc/EJp0Q79PUtRl1WLiIgCfVP9OL38hlsBicUXIDa8mLngpibhh6lNkc
iAJP3TILQCEGJcU6Di0Zvb+y7UTxIVyGjNnNnxWlkNHpeWOfFjcApy8p3JRifSTTz6fXqDy/pc0y
iYErIZpTh19mhP2ZyjYE+vORKLOJ4eWlorwvP43T5VTYc2byRB7BYzIlwBh7e0FmAmh9nld51N5l
wuAloOWsWGFuXwevcXCUNmqkv+HOHo7vMt8ChkAVwbPOF5m8Sm4VxM9dUOr7RVlyH5hhJ3zPV1OS
UbbfFyP1+jzly4ZQX+2dCzc0sFIxkzQ04MgqW/QFLMmlZz754pjgGW2w8EXpcyHV+0uqshePzRQg
ylT6BaJtxkK5cS7pKZOePry1DGnj5CuVDd0MBwwk/7o+KFCwvY2uA6b8Of8G26BPXVK8gkYZhDPM
64p7dsBzPZ63RAdgJ9jXcuw9tXAOLxu3TOKS26PztjcLvccbYJl5v8zDSGl2bef4Fgqvu5oSkSKr
cXXXfjdsyuTb/5OD2wR02oEOAWRm1+2cgpASHOaVaSuumJnTpj8v7z8UMJcCJbuK+yUi015VBstw
D3cXpF9cvZ6TTa26R7j21mdvU+BuGwyKZVTlebY+LBtqK64ui79R3D9VfIUQ9yNycI82L553Hljh
GeiVlGwQVK9sJYWc7KoR6whhkG4uJq+Mky7HaVbVle5so0ItQbH/I9wfdC6zOJ64svOYVtfkEki6
Hy2U0O8/f1wAi7ndTWG8dN5ut3o321VT4wTDEoUamnheIbZYSawYjmuK9LDOd1OLuCkPO+9y0RsN
UK42s2/NcQUqM6LgvrByEQfHk3s3WuDtAz+FY6w0hmvcalGi6k4HN+T26EsiDAIh6wdOTgYX3JL7
1W29sXD1+oQqi1Md/HKDNwZHqy3+fwP3MYXXyRM1JomuJl+0aOuKwhVSew8FsaXs38iBpRHMOQXx
ha8eEcuAr+J3N+LvPNhGOAlr9HUjX+x6SWOOj9HS+QEn7XD5Z0VE6G+eSxxB5gQgKI5mHXmYl8Ti
4ypd2XELyfMmACAxRrIDKkZtONup/p6oXlKe0sBWc95NFQL7QFz36ZjvEdgIus75AKs3C3LWqK91
FIJBEQznq8IJBB4W8A/Lx+ljPtmBcLt2ZYs94HqYHmKg/F2B1gTNX1VarvSSRN0mqSEA4agM1Wo1
/OGU6Kqm813t8A0AozFA7DLa9PY/NMm1r649QhIEz9PFJxB8fnmivXr48BpueruV8yNFAeb8tTqF
uh5zvpRjPS8oXTd60YAPelc/lUbnqKdHyihYZlDe+uDb4smB6/zpnvrvNoG2l+7H9kJrQ2kNVBNW
zUsDuRt+bpD9wAR6sXexIEzPZQM5/wLWOjnES7K63AmjJuTIvHc25EJa/LQ/QFwPXBg2eUSSkclG
EE5sH/SP8hxkcoOKDAi51hc9FeZeATbaKQBsP2M+mbXPdsBOlpbUnJIRpDK4TCstI/MhBynn3b5C
YgY2iuICPVwPvI52IXlBWs0cEpc61ji6nleBsf4nEbr4NHd7DqCGLRbv1pxKiB1eZO1KF0DAJs9K
OmQTo0CoZYGBy0p7NNfMh1Jg3fKwVMzOwrROXqG2faGGWRBBUO3oIctaZ9MLBNo1c/vRgkoJNnd3
PsrEsbgEXgmFSCVmtqJcRuapv7AF6QegcoD17+tmJWimJ7QCegKNJ23KWP5NKzTiD4jDzVhewNOf
YaPqJqH+7m815gMM92HNKbOzc/Jn11oj3P4HSdGZpw6WU6FORIoEpZdrNPQ1sJi5U2dNQ9gTpR8P
iVUtG+wIDJN3D0rNyGNvQb6qnjim438OKaIWpsQvXIxlNxutyBKH1SNXpeHM6TtzaVLZsj2d4+H+
vhJYEcmTAUA2OHjwCr+Kp7gvk/uqZOUUcr23nldeLcxwK6aJzSsGhYnVVoH+C0LW7oeGfHt1oojZ
kMhj1J79K+ugSFXjaneLgGM2pDohmgJigB5ScOAxhk2UrTVyRN6tQ6nL7TDG+vq+tcHcrE6O8zoF
XjSQ5kMQtkaJGh7itKEGwzG71w/R75b8+XlTheu2dTcggnVIRr8cilPTmaZp9jqaUkcNLYmanAdb
MVr8nZTqddU3Zp+cKlbvSxfOdgzLJIg2HBUouzqiKUdMyg6+Y2vecDaTg9U1ZB5hCwPixCoE1tyX
BQpbfy6HLjetibSFzdvrZitKa5Nhhqo4EYAVMbg4m/7cRbUlOhFcGjrkxRu3tdkZau9zQz9zSjQ7
aaeZiuYhjltWQTmT/pE2/QCRxUODNlSMA7ARc5vfZIkL68OYcaiR0hPPIn/qXpZPdvgyjyiEOg2i
RGM4/2lLaJiZqSV9Ojc3qnje2vItKyAKp4/bVbBM3jQvMX3jXQvFZQ4GRFVunu+FxwPz4fC3rn/3
45dJOHIkQT9Hk8RKvse2ZYv+gZ/U8Of8lAnexz6D3yY6D5PgC6Y3Amxrr4vVgGXpI0PQ/JZWvIIA
T0s0Rmm2xbKTR8uDEaf9cs40GWf6MxX651GPW0D5i5q8BCBYtizvBRt/R30UWoiZq+jdHcIHodRU
2fAP2c2NgcGI8atYbM8dx4xiExwtBTTAuPRpAAZb27g4aMMh1oPu9pfcMEkDYG4KJRz/+cyDq1QC
g1w+dcsE1S0YLzk9NsRu61fKvdNk//as1K221baHGRXWZU/jTp1lnKGq42QR/OrWk0LNU+w1GsVs
CBCHlv2Bs9yd07p34X2ST4QbLhvOBgSBBW2r3B1ptIh4CbN1HAr6awBvFSujvNZdxG4a00vZ5MdE
2zSEm/sY0vQ3DgDqwz+epPqiKioGQiwt2cbeJglk+aG+7z3U/phbViZwaZNTKRL8nF0WAG9g46Le
Kh6BuEIARp576hwhdVsSsn/6ruU1rpY3jPMnVCEi6+sYtYXawBMsKvH3N50cQnHoaA0il7XD+iz/
GAz5gDWorVRJzdZPW/kU9Q6JBLIvmPJuzsyy1sQhhc1ER1WhGcfAVY1+ealXYbpGDzUTLxlyU0/l
03Twlj/FAekl8xVA2IgjzqrMdnZxSyvAeJrpHodTvCBV/C56YmQkBEDsm2IfBlJ1x/PrWUmdjACd
Oyk4lFYi2QkclfHsO96VSHmb8O2dUpDqcdS7Uj2u+Ip18fbrVX4Y9f+JNBV8E+auDYb5tSVXTrT0
QBIhjLx7we6DoqT6mX42pHEQkbhEszhJ9q+LowpCfB7AJCtYmA2WUFrJHCG2w7LXeee3ZGcmkJZW
M6geuhNfvMZwbr/rdJs8XN4g6GJs+P8T/0Ywe1LwmrWHva4ns4RZLFwQOVg4VDQnmFRHecxBhEo2
6qFYCmLi1jfrTUSPqcKlr4ZBCLV91uPCDb2o5ayQlX7yLdTVL+XVNDkBugOawplrPwZUDKRjdybN
BoIEo+XY72C1YATkrYSQGxhQp6z1+uS3/l07bK76VmPWzin52bw6O1C3LOIU7tbN0sfqLktdChqV
FnYmMZuL5C1/L7Cz1U7GVoN0hrNS3XRNl5J3/NVQqeg5RXQHCfCCYS5TM3T6VZfkh30y4u1smTVz
UqcOzd5IwUeFCZp9/BFz0rHznb5bEtXPzr/RpbN5VwUZar4mtFwP4llrCBzAhgxcP+WtN+2kCIVL
dJTLwHpgzHASw4I2D6zCRag+tTbI7AGbgZiFTekB6u7MGYKYCb2QjYe8qZX75Uywo4SclVGHOIkC
tdT2PWb+Sxxv9ZpifEZ1N+Vym2y/mANSelm/aqJBUsTfwd6nl/5Uh0/EkNoCSMsaxw8GcYmqwKrB
+oKT99j10rgnrtKrd1wDphjTuzGWT8PcxeubnzTa0T2PvyzM7/oDLXXWZy/92Z1H+qd/Y2bApqIy
fWZMqxJQk+rbbjnDFUX1fvegSLHTIIVK4nPpM1sjZjUOXB9XC5SGeYaZ8AcYWzGMkHdSnD3pZhgZ
iL1EeV8cSnAFSqgVwiKfKN+yUW1poKSrFrp+YMMmpovbhgFC/x+mJAhOWEEaDJvHxypSBoOmExSW
IETw2JXr9INF834zlVux6kpKlqGEQWPRa3ZrsYjk2OYSZ0yutBLLVYA+5hcT9tWzlmvHrqHuhDu/
WIG8UdNS1CZFvuXO/fORczINwUyOZWzcE0LHnX5Xm8GRfHmwpr4YGVH0IJoHl/+HpiUZ5r+YqpRy
MbhOis+VmfQu3CKZ27OhbKqAF8RpdMLEMFyJ4GDRDnUNVPQbaQpEQUXRtpv83IQz2hcktKCjxEKG
LG78MjqBCKhfeFnhteDerPPe0UbZtw91EUYxnNySo4OkI+Xp/kp2T0l5L1UrMigk7ftu0zdLxy2m
+Ckx17X+MLL7kMtdxTGzjPjGNRBkWwwfJIdkllXUpWN8PUgY+WILBp6QMbI04jCS3SN7WOv4sEih
UIAyo+GAd1aKF0raThXMoO5gZQAMcpGdF9qQkO86sBesKVVXKTqZtH92KiMImAIsdJSb/BngtLNw
dj1oSWrXw29Ayjv4ytE64O+XJRev4Nl3yXgJ3/b9CfpisLwjL18jZ1I3BxdFyQkBVabd58L0AA4o
J2TbMC2s6S8VJzFenTPPP6SLNaNZ+pZ+LuL6AaAuZT/E2zNxamqmnbEK7jJGed4JzbINyL0Hidzx
Co1XcXkQntJnqLNPnRPjzV9ZWhgciGSep8RzgZLQu7f6hfm8TxvOIUxNy/dEti3H6qi/R5Dh2E/l
ffOTl9tSp+2hbQotV8TEfHKrO9sbuJV2PwLg7drFbcMBQGv70pIiVc1M9reeK95Y9EwoRyOn7nKx
CAo0uw7Vkz5GntN354Srp3k7iAScbeazFNSdBnLwA/N3qt1dAdZSUHv99NNW3rJdXbZEo5TLkJSM
tqA6FvkyXyz19svRdN82k5Rg2nyvnpVMkKQBQpdLhKD1+T76SNRwjG8s8xv7d+qJAT0uWAMYARv7
JzTndeF8ir32fLXUZ7DWvVJMWUaQlkJn/08KLdO6km5XBTqMD5+6P8HGXihDvxlQozH4WcuJFmr6
8uTWalzeTp2vYcqiLf4zGTS5C55NMzczZOHr/Im1vr6AzGb1Y2oUHpWlILwg6RfgyEhzIxKAjf3t
swrhqHHMOsxzu/3ul7v6EVGbPrKdbAnxH9Qs7jM6nZLy312MlwP1xFrXjafShBxKbAKWVpiIDrqP
ZlJezT6Vz5V8q9vD5y8rsPiH+RgGTuoLPPjYf0pVD5uxhgGA6Q5yXcDn9JapZWY2fGtiG3OkwhWy
C7YJq4crT2U9wasJgUvrokIK97mdV+Taj3xdBrRgKy8xUBdVLiKzLAQiW9Vcbmw0IMyBVF400VTH
DShWGS2BW2l8gySnBMI2nNDwhPpHRGWI1suH9JMpnhePEKlWFgry8BNjxPCiR2PkXCwJBgLBEZrh
cmb9MBqMGadONBy6b8hsODeDWTj+8D9pmZx2GwoXeSdFHlbj9U8VRRTLJAOm4g+RI9g3li4PzpEo
Z9AUlfqxn5qeyCnAvL+kYdTAIifBBun8FFoWGKc5CIkf1iNeabBg//ygW+o0cNk+q4/MEKEspRr9
S5+0393bc3dnmTJ2oYjAHIved74JcLcAgvH1E5foOdbUzeuyVbNI4C1ZGdurNFd1cLfN/Mr3c4cw
2HBWOnX4i60ZzzxjVqTEwzygPRwvsfYTrh0qoTT5PssLvuXCW13jlU7PJ7g7molhOM4PXOx8f8lV
lJuxt2UTJcn1za2MOLaVJ3jJ9PAPg6t8l9oq1v+MzFa/AHK/VmsxogBdVIgxlUyD7RNR4fPQ4jzm
+FY9jv+CT2Fq0k8oTLLPIrj9cVrZ8A7uR+A5HV7dwrp5hqwG3Ye55hZlimkmtE8Sa5uXOrJ1SxZG
OFFi4pPVyYnJ+WRFW/a9SlqXqa9t8392laGRvT2ZLnTwwldfeEDdMubFe2M/MaZcGRCDvs7oWR5k
HZjnTciUstKPnTzj77uzXCH454eovsEfZ6VRqwy50uHI4bnlz8gIyE58O4pGLZJVYf3YbAJ8Wrg9
JbrzYVk+5CPa9SgWFLNg6r3qRjkbMyhU2bvaH7VcTRGW7Vbjel6PjYdK7a5tzyF+63f0Ylv8EZOr
CrHOmy4rPci8nTVc85ptKnfOf6fPReOAFn6zwHVrbKChgeirLY5sQLi56OfIAexfyBliAGGJmOxZ
b0n/AKnyXbv1whysOQFTWsi8eJDqm1s1Cu/WddjSzMxMt+bamxWNiCJuxh3p+lEVtGS220ZBTsNf
b6drvPpl3aSpG9kWyY9tmjs3IvYxzbxcimYTXZmsjVUTt6SD7nDKAndQwAJVeZ9EWTHV5r2GeSzM
qP452pp94UD7QqeojA5Onw4LX4DO3T4OVuL5j25r4q+yEZE/fcOFWbChAdHZ3jXXPEuOU7zCMgbS
KbHqON1F6aMYuwod+SrB99p1SrvF8uDvHRI48jBP++V3RgM7a4K3OIo4eeIkDJgbkjW0bftD3bA8
gxUEu4KV8kDIW71sIaUvM+WxO1mUxbQuireIXTVC7ENtl7AiZnPAptaQKk6WWi+TM9E6bZh/UxoY
hxmR2M8Zf5RU0w2s3nWe0ZE3woRGUAODv0xqIUpgE6MJHc+mtAzCf6nBThDXo5TJliZQsjR4xrLh
3xftZ29PkyUdtCia1Og8K+3EG1enzC1avNL0+9ucMM4iE8Rz2GEfMID1xf0g579YZsyekXYHpRLb
1Te//2aHPLgEfp1yYeerBnA1tkKGeHhhvsi8JpL9XSDrlxkU2vrK5/Uk56O2FUz0b851KxmPj32S
DcCmqVcH40BzOyZKgASiiLSwiNINlR8kg6mHQ+CevsTiiD/x2i96YN9rhmDHLC4Ke6sI650UMLqM
CuR37bqLakwS258MwCvkPH5sH7osKkirv+0+KY7iiN2E39cXqcn/+dKFOIi+6mqgPLfibq7zOUzs
+KZrpE/TG4dsBahSE6T6kJTz3EHIpfOgX/89gVJE5M/YuF93PPFn7kaRqSLe827wqjUitk0lhzTv
1tZI/0U4HI8xPgNhDKB0oH38hfFEo4THLZ9uqC45Lvm9GEkGmQKvBHFj2apQquo+QSwDOwXmRzsI
NGAeQRuCdkSUe104Am40+GGPkHlmWGAmi0+THwsokCe/EkDavJBV8clYPtsLDfkp2JPr4MZj6gGo
qTLsRQIK2v4QgXZ1L96+lIUwpKUiTKfgKL7OuDw9p+y+fAPe0WrpNuXy5UlI9QBffVBw6pJIb0dL
awoyHcS3p2J8fToEUnxlLUfxPOqVUYkgfjmsqLlI4EXtk5TjPSsUnhPTQGlFqsUlzw+MuT2jYv9G
dhob0Uae9Kt6xHvxQxt+6JbU01qtspMGHNhnHx3Z4C/jypGbNkzDEC3JGdM6uMuovU71Ptv7SLp/
yKcz/p59Qy13LOzNh9wnvZ1L+mh/m3DJ6GXS1v/Z+t21ZAimuuFwmsQ+TaMvHTGEgLM0qD1LbGUH
nOEMa4r9MhS+nJi+rwPX43GLo1eU/Pe0vwxOhQrnew0hKEV18Hy042C36mH0mMjfZwyjanT9PE+A
gfVzQ1yjxlZW8SOGKUuenWmwNFUevNdjBa1l0aJvy6SJ0FtL1YPfhciTf9uSa/xThVqokQtzHmrY
tMgiZ3VQxZ9D9OBydefaCzZZJ8yEgzTKJiE+bPYTM7fzXwZb5q9eSDSiRu8qkRfkh99KbsHVnkAp
cR3SgvsrxIdVqmfwWVv4vXcqPPs3PUmkzkaRiD8g3XUWK2YHib1LD1XWLffPiAY+48hPO72NfBt/
fGm0o3yMwnpB2cyycvhfM/Xr4P2UX8Zw43uzWYEDPQ7FosxKAOHn8lnuXZ45RJeBlhBCof2PAGf6
pPZ6IHym/aMyyrBi8mpw/IxuBkyOtiFnypcJFLJPZRXriaF8Mm//kStGdMDsuXMSUd11jFGXlWO8
hGfsCsdOLtn+4q7C197Mi1bm3bOvYq4rO1hySornMtRcM/inrZA3ilBvtBH72MEPAfa8r8D3s86Q
9VNzERWY6A/yi7JWBn2T8RBwBdP5wniC5gJETxfgGR1ptr2Yq73OX3qlNbyljw4Sjc5mXncwvkT6
Jt317k7S3iVF6JttLwxpzQtrVyNs244X/Am5HDG3zi72il9Lb+rbhqObDHozrLAmOFlC5gdizhyI
VIbJ/sewaN5RuZfvNg8IHaA0S+e7RvO7fUjEkN2TBEn3mZp1tfJQQJNujCabh2S3UaqJp3XwPEfU
vZl2Gs3rVFqwg2yOEmDxt4T82VU1EYVouCtQ7xqLXjcfIvh2Ya0gFUUaZdNi7R4dSgPmrqO6yN36
g0r/sQcr+l6NXqQegXpditQf0InTFMwy/mq0gGF6PDoTTlHy5ddSMlRCCVvDxNqT7ENlVK+2/byQ
6nEizHcsZJ+VY/NZL7G7jCmHzvAAne5YhgbiQzJx3Egj8R2P2v4zIAXeJxxThO5gfMTEW9Uwmh99
0tiW0cLPfE/yi1sxEEUdVjg8DkPrTupWGicAQjD3DhcxQx9h8lIFOMhENDvGEaYb2b0LyL8AnRex
0oR8lTLSEtVYeWZs3rifSOy+QXG6V0r5GFQOA697rVu+KreVehQX6531w9S5nGrABVyx4lBfoZG+
nhEnaJ54QoSV9Z0yhRdSHNol7GF2HvfCsXZ7PKTL9gXBRe316No7q5Wl1vLnZXVqsAb+JWEa8D0F
JGSuNm1OWGX4CevQBCd/w+bm+9onk6htZpXEDkNRmVdT/84I5lbDiEzVb0f3tlOdHoSaHrOnLwpZ
ZTnezq023Gu15pp/DMS+cTf/9YcFapboRahgvjOX7rKVsWnkQDFjdKCWsHNJrdfhgnarLa75RVW4
JlYCkyOGkxyxj7eNXr+qxFxZv/AR6NhusqBd+yP2DudB1IdgOqEIxWcPyjj/+D/7Com8Ju/fdRjQ
cBdJU6V3Y3TfYUyDk+0LGXAW5TKJIheH7vy0PVoDkWl1wdFs/ICeIgwBqMPkp3rlQWOeSnLQ8c9k
aVxDVD1Q0uW0Rsf/nCmeSJjIMwvTEJcLymm5nsr16nNbrVksAM4zwp8kjQ2Fy27xhCaaKYkva2fk
W1vVcmxaCDw+JeIZpSbWF6lCnfP9oN0HyBxzvvDf82mhOjsgrvV+zk2A+8zjKgewUC8JC8fR8Qj2
Z2dlx+3doLAjCuCFsxWJc9FBGMopdIjP0ZQ7Cl0IpGkbQaab07FAl+uoho+kEk++rHFPUMNqpYfA
Tl7zzJOi+kKth5PAPWv9wfkvTH3d2+jtdFmutjUoPTVk8omzbWVLQ1Vqy4s3MrV69M36x1VQ6e3e
29b4Y/ZfsHCDgjGpCTLlBxMXkAcX2PjECfkSCI1qkP5BIuTCfSE0z7EMRryPscQcD+v+PKPTXC24
Ie9D1wROjjHyqa/hBXh0by3yLP6AMJ5tNl9GyLDiOLMZ7coFwZdJ0BuXhEALEfT0+R/ZF9EyZcMy
C8/DhVFIKg+1e50BB+5Lye1MnN11hq7Kxd9mLax2tNmmsdhArcrTjVbch9+XNohnxwYvsPx40ePP
fZqSw3Ck7bjLW7/qGksDxbmvr5FOie3MXHCwyhfB+KZzyMh1U6Zleni5KAi2bjC//P2dvYfyaCrA
BPJQNYrKS1VK3r+5nWcPxYMlkTGB1jyzRipsPMCbPWWWkrnb3ij2V/u5crKSh/GdMdg4lsb7sb+W
LkZkBSA5hWMnk7S2vMgdHmdWPT3uvsoHyEaG084k3P+RSsAY/JEgGEGJSNmqSofZFumv69RRtEwx
OjDUsJ24AiMeUhEL/pmFBwkJQwVCzH/RIka06zaiS7j1OXjDPBIvtxFmIP9YrHlYMADRO1QmOONB
NpjdYVZQpz+OE/RUFk4BNmIyJjm+q6N9iLBoFIurkBcHH2dqPCF4PMQ0uNHMOOzHW2ZnUgunWKcj
PoVhDbw/+7Mh8/SikcyJxCr7EbwPJ6aF75qArOasSlKVlWil3Ls494iQ9bFdmLDOER4yJxONwAW2
pwXXEc7CyuCUQVjSDGkArBLZ1tWPTleoCEVfaxYfC+4fBs86zIKDOLKli1wYMN1/dNb4GBxcYhIE
buZnIJOTj73dVpWFZiFRHq9mMC7k+S9/TwhRvj/SrYTPIMqRraMP4dPdYg8RG5R+QqAn7X0Z75X9
IlFcXlrFkr8zkzHQZSZ/qtUPu1mn2mt8MqIe2xWy4EIngrsEvW1Y9EZCaPafZzzUwckT2S+YOPi/
kaF+B1QiwOciAZyjVDy/cFoOv3Z3vh6ZzB4iGoTIvtAU6rDKEiMPvNUZ+a8HnEJdbWNbYshfNR5g
eJO4oV+wmuPQ1H1hKZyN5rL75k88lzSEH6R7n8FNP8mM0N0piPLOh0+Vjn+YRCVYO+pDMZiOQ3/f
TjLHFVSE1uRdmfH6QpAz/D7z6bKyJcu3ZGRem98/4k9GdwdEC8nOxf58mUzZSkhdX9AT5oV0DCMU
7xFDCrttDkaMMmmwOnrvyHbTvmkzEMk1VBs7CB8B+t6jaQH7l6aJNQMxHrAtGJioIptwr8tfN5M8
NUE107Asc6RFNQtkFIScbTA4VBGBOvkvR5FTJ9vmTGmO/WlNLjEyUWM2TM2nsdROtLLCaEy0a0dz
+TRgOM6Z9IO0QCSZpyKeeZV8/EkyH46KSUcxJXh4kB42dRTR1t72lbpHdn0hMqCiqM7XamDC4p41
yWDlo8nZApW6PV9b7CCJsDyNq9KUU4PhFHz2+wi4iOW2V+dwfOkhmvxpSkj821LNBHBgiQPRQT5c
SCv8RN/izzqivMGjcV9uvwlBZIUpMGl+hYBhGpZprMpPEAcNOZJ/Af1tk1+F9d9zFkFipF7ueg2F
K8aTZC9HF5+XnsTsN2MHRuIVORFSalB8gLUoNqfvZ/z+eTR5ZVPYyfLsyc53l5j9f1Hfc+ixYkUG
Y3ZzZcdV5dzh+iUhhi7pmXevjRq9p/itciEvvGTa17xheeB80zhH8EI03arl8FXJcflEJy03qrYV
KFF8djyDw5ygjzvhcnwqPMuWPMIVg0LMq4ZhonsBY2b5HHWwpy1w3LylfBVSuC1kf3UUF/QFAOb1
J9eh0HgimJdFpZgzK8mC8AFAP+kF7Nh6yyKO/T+po4+g5qUaqY1MpIhM/A26IqFbzikJ/Zq1ibNc
NJ8JpJlj+wheYPfO49q1Eco5fjRKoCvYy9dnuW48FDPdTH1naSeql3BUFHRr8bQ1nC39gAokhppe
cbjUdz1QXbGe1ZYZF7wLE+pdUD4Y8qBssZtKUUW14Kz7+nEcQXNB16JbMNt/ra5Q/wnL9EZfQwqm
1qPfA2AttAVtom//AvdIm/UTwWyhKh9m+gBZ2AfQb6BnX0Bb4XVXkxcFnQbYCWO76VZPiDl5a+GB
5XQMSRiRou2algvlPw0bDUrb6G/hhY4wsX78/xerjGaxIxu3q3xDR2XJ0uqrqhDgC3n1imQtVfQn
92xs+wd7NjBxSfKpuPimBSTjveeTxSkbNgVPfNknAhPccHR/wPaOqrW2DS6ClAnF9ergveQq/2cB
ibu0xrDWzFe3hagRnUFfsJUvNTsxUj3SlZb+KVjoGk7wh2r/cm/gFibRlW5je/loUKgziDNNjGrf
u1AOqv9nrj0shcPggTWQA1kMQDCEjYnAqaVFXEYP6mgZybIIWRM2b28OL8pW6ZVN8dm0RB7xkG9s
hEVbN5WuoINLPQulqHP6hFuWxrJ92+v3MZOWHbo2k4eN3Ay6s6qKKFF1whfbTQNa0cEaGpFHdLjL
eQCvP+E4NNxN6p0MInHQU+O6Gmz3KdRDcbG0Vg3BMHgEsjfQBhrDucoYjiqZ+THUCmBywCqhB9Dt
Xk5Vf/FO6V+53dcVGIXqgLNfTD7kc+k9Fk0/5s7iE1i3QnYL/1Xc7mLp4TL0NIqf2pL10VuY+AkP
O76TJTh106uGYl7vqZyWuCV+Y7s17HEAbpUL4efa74gKRa2r/7AL4dGhWkO4MHUb0f7V/wqhhEYF
NR9kl+xE+3s8B4nfCDTl65nnovdrGU8QNCaV9hxwgYewYZXRmhgPQCnQ4++0N85GLytzYml/joGb
Tk0Uu0IcXml+DUTl6zmev/asnaB+60Q4zeYK3ST8IyXaqaC/X5XQj83aoMZmXEDynYgaidD3wf/D
nu/T8/4CRnXyD4lbQlhWdWGUnmkiIlSCcdvIGAqlWrPh3/IOGjqlDC6Nd+6ksxHPZ2ygBYgkVDgC
zXqFOzPZvswfW6EGTWChXSmZIEMmGTsggazleGwJaoo2mKqg1+1tVqLRTBLu3MpjqRO1YNoBxEwR
bJVneDppJkULeDRvsChSEbHZ+76NFs2EMWHpscttC6WBGU89w4fdMAW83QGLDFXXvnS9DuXFgLds
HphUks7SVSvRYHrY45Mb9vz4esi7o3w2EpjmMuSJUDVW+ykJ/diFx1lxPMfCI7NjDt1y0Yv8nx6f
Bh+6jOdn1ga+r3QbCyhW3cY8cEDYrcYcIZ+1enn9W3h67VCsJW0zS4t1TU4WTZc4A8P0sYnUlfjc
FzcGNE2wtNM+std6QVFXVG59ynlnZ2m8Uqr1JAbqGkJefu+dP2EvR9PNiaI2nnSkTw70Mjo4R4cS
jodBlC+sqo7uxen7oYtG69ASrPQsIsGBRwRJvkdfEhHAU57vuSMcb6qIlyhFOoHwRgHs6vZ4r5cv
6GOW281tC820z7LJ7za8FQ0dt8p8vFguda5Hr7kYODxRYODWZWHuLGwhAagrmMGCeBlW7LFfP0n7
qivmq9xAti1aWG6qBSD04egL+0zVZ8Fphfbnll/T60KTT/rTidT4OBLv/78NgRnssb4wiFxrwByM
i3JI3Y3uLH59zxTDP0UvQ4H2DAEhQc93yIbb+7sek5ornFsWijDS53ee4VOynZ1ooxtkFjAZK5Zc
0Nx+fod/n50eDr/u34ELT/yIhUkQkUC7Y5pgsSQwyPoVP4oEk025qQu+fpP/g8bZP27H38s38Zsq
I6L6owzWAGp9P/xj2YMITcY4M9dDascmKCx9AXEfzQjEmhFXptsTB4c+HZon6zefv1aH/BBezRU1
G4eQSiWB3pqbxlLsE3wAlhYTVISKIBow0/QHkbI2VssD4Lap8vmf+6h95Zn/hXAIitXL7ll/lYmm
ES8pcgemIefJLZzf0QioUcYgonJ1mCVohR46whujZqCzjEkndJX/bRBZJ+/Fg29oxaBy59icMVDC
2oG0JVT0nR1r0RDXO/ETgCFriN6efBIJC/ull0ZTsXQIL8NkIfzpa0fWknD4i1AT9puQC17pB74V
Jxc700+YH+9epy8Wo/YDkcMa4XhyE905NTbLDijh7kLVW4QL1OdqfyqkdxWrR4ZzKoeLd/fVbN+v
hllqtUoHkEDp1U4sFwKnXelG8Gk3c3zqGYwbBhKH+0QWZpkPlMoRZpDE/QaFG8OVYjT3RBjiOKyk
grhyqM6aJeJQYJPbAGw6STe4GGRjT8EADnccgQ5hxjNihvMztaCs2cmL4lDjEQGAc9xcyU7BfSOJ
cXx6P6RSug/zgiHM5hdI/FPl9Gvexg1+Pn+5sje3/PzULqBIlc1Lo5IfsWEbbfEvW4joIprWd1Ic
Il8Enj3u/PjZvK4E4/vkVeE0K0vUZYithBKlmByGsx+xXFPgLkIAg+1eq72XHtmRUrDMOuC/qnWn
gmcTxnbxskOmfUeukl95yzoNdQL1/v8zCQ8pzUOdzKRwX6IBjZid6JH5DwhSCjlw3tckvINnqy8R
yGOzNjdA+YpHY+krpYvoFmbgVHEcI4cUa9L2yvwcMa5Gkjuqog7BHMDPLlrCFUTsI9G8MEveRcce
e/9pHm7/y0M+tQBQwV5iKch7ILAP4XPmt7Bu/FuLhJq6k0COXg+lXEZhb0ccfObT9nJk0IDsEWfv
y0Hf4JPGhglb0cxrFew6RUhafpO1llZFPEWRuCXMAMl+St5p6q/jvkU0ra7KWyWTOjHAhg0VESYL
HdjISw0wI70Fus9nCYiESV0rifX2yly7scewe6TFivzCEtstYB68eou42k9N7z28jaNYgGl9Rqi5
Cq7LMBxGt/vZK8HOTuAy43AllvsYwO9uGjEh1Dgf/F7XyrneOg/Oiem80CSzqbD0Y5RqbUl9CvDX
iV+u/fh6XwJnEVyCB4zyYSJ28ygXM7YxuCpL9uqfGoRoG5Q+rHN3dkQgDQ9hy/L3JScREu9iQ14D
m3mauSW7aglZGisbgGEuaa4qSDD7qm4DJwWhA5lIXmEksFIUU0x1qbGaSM0T4QecKFRMdRyXdySs
OwMfOI2oVEvbGqET/U1rWHiwpY/J4f8PEnQWbeOlmFt7S4v5/Nt+Vjegrr1lqN+Rr1FvpMdzfRYl
a8EsVPiovZ4a2wCorVCS+C4/fpGcNy0RdwLM5uZd5natXSKQIKXq+qP2hsL/Ls1SN1RsarUfhTlW
uaOtzYcRtqe1SiSI/AKHfvgWZBrDrhp3I5ffXsJQaXhlgulmFyqVw+d49/xqqIETULvSaS1sR23G
JRXezNvJMdtVA3l5LWayry3M5/tA/fA65dIBVTgRIUbi09/fOFHYVd0JgP28wPkPGZe7Jv2ahDpi
yzCFoeHcs4vY9X2rZCJckILM9jvOuc4JTQdltJr8YWjZnDcP/wghOupQwva1+CfOYDDn71w+IAtK
adnsA8xIcTIpSMBzWfe24Mw6i6xCx0LZEdPWHpHPKwHrOvMGON18bbz3OpyUKQO5eKsf3K8bxq4T
R1mGPq9Pi0MfsFvXUn266t+Vf/38uUBKJvhKwTEifGOZ7nNBWzsGo7s/jukpp9L8+McV2PHxXDNH
3IMCy3iUAhwf3PWtgWN8dcj0FFcvMaIrqtyH4VAyrFGlPg1hSdIdSvA1EF5LdnPyc9GRtEnKGqPD
L68LxAkv6WMJa7TdHPuQveGqC0jxGEUDVkg++49y/xjjHJpbZxzmXeXSbz3HIlWr6QcKR3P3b3lj
x23dpO3g2EvwiUHwh5/wbNEJaFPaIBBxQkE1vvat7L34TLCUuD149vn/SfEAP6vZlUCdiKZQlwzy
zlVI8uJqN18+rGIrFuC5AQtAjqoCbfh8OANI/htAZTQ10Nmj5p0DXff862CsAU0y0tKxw8u8b6TC
UQBzOrbniV8KHd5egP1hen8hrZKGUtny1NBF9Q4C2szAMq5JGWyflul5XRsP0OwMGItFiWPAX/Gz
57Q7ExnbuqO6FRWq+pAZSaWViW7Oi19Fs+/m8wmEpDd14R5IQPO/G+zzeoTZ8cPuayJ4zSGMzlQh
lnUT1qKLnMIBQuAHsJy/o692d4x0BwM9+VJGxLCyAGlUoLCEWspyTIWTMleeJXTxGRLhjwI3KRL+
2fMUvaTtLOwcdASFVRGGxaSqyQtGrnApjjTqQ3kmLOdJfsADP4sn/yzQiHUQEYcAp1KX17oaWpur
0CHQLbPBFgw6UooeILqKDBopSOfgJa7a5I9QPqnKm6e2ALESjQ1XR5t3BZveQ5ZKXMLZmQU8Xl2Q
KZBO0e2h+nidpISiQkEQSjg7IeOWFopnY619e8HDhm29FLz3+Taz9eFuI3Bsr4Zq8uxjf8vZzKkZ
lPi6vpzbr2OUwcJtoazf021DGVkjHRTPFFbEgVYFRs0DmNxmfaf8JsKXyrKI2GPiK+yDfPcOpmzs
7Ligydc8K96ocYQwFu30G40FQpzyyDjv/dtI/8LpbUql+uYCpfjjKTlBcTWkBAl0PhwCrEKqitGe
f1ga508t6h4zMzhWAhTnU71odMlRDyNlHChwxVIJcrJm5g06DyIcbX8IPALCz2DRtRzFVSYAEZQu
WJVr9dzVcUdhr5/oZoH2Iq/YgvWm1gp4xok1t87X+FCT+9ofDRknh0YQcMjXIyImv7pp5cMg+M3g
lPKF3wJ86xOFl4qehmirdmRoCMXjxJCx8C6govhy4BzZfDUFoaw3MtwGl7l1xPVGwLyYt6F/jPBo
gf7qDIkf1F4TDDIlELDhzLTf4dQ/V+zwI3lj2qKhj7lJ8UHrI9yJT1FZEgo6H/D+llgxW1Fkn4S3
h41ST8DerW4uz0NeCEFERcFC1+3Cj/YTKlaN50Bhm1XuiPuvsIOZQldQVvaRY1oRmTDRnJNnTjha
0SmT33lbB5ERbWqZXjjuqw6+kY1rZITw5Rmoc+gvvnFie1JqoDqheCSbD5+Xi/2KxfTDX32j++y1
9mLejq0wIiDHD6n38m0MFcBPTGlsjUTAYE7K/vgT0vgeKTpk0MqcoGbaKIi+ii7JuJAjP+QNtchH
ogbSe3898VWzYTf6TEYgeZUPkJEyH9xbXF0sQr4Gdh39kOlYi1bNaeISNvDejC+aTXL1AzDaXZ9P
VoYgQkOqFHsiSj00xdXvD9KRlcQLykG5ZBOaAIaLWZvBmj0ur6P49vObWB0999Ity/pcqQiXH6we
dWQH3TYTa/rp10fOJjBwAahkYJLpovtTon7JT5F1QRW5RdSgMeg6UI8/fvr+APNRFU+e9JuM2JK0
jlBGFxXo1suf3FxRYzIaBMp+Vf5DajFgbI6zQGQv6NfzYl7ZylIRmiwp5jwZdfS7WmYc3Q3+WaRG
a/MI1AxWjyEoWzKlT4dreAixZsx0DNxbkmPXIo2JDDctL6UgDKWzqnAMhm8cCwjw6KDQxVzcXh3L
7vu3kEM9lGMn0V0OUkmLj5KXiZ+93/nkbVu4ZF+otN/OulKhq494TQ6gajOODM48hnr2D8wOYfmB
NmEwCiyaQCqNnGDBOCeQwMQBw+YJ9V5r0TD2BM6G/BlL9mJumNrfjF4R8ITXkNtvtCOjxJCrL4s4
G8MeWnKudZTOTmKO2ZZnytmS9sNLsnraHG8Kos2OM/+/C4CbMAal0rzuVo/EP7E2RTixWrH1/gK9
H8xX+H4LMWsCQ5jx/iXkBCxStu3yZhL5Th2hW9HV+xIo8/uX1JqsLOURP9vVSE+v9jX6YMwfX7yQ
C35c0W//m3g8QqBUQUTEDqozOgVaYPDPMkgO0+m6XGmv7wmA2LzqfydYHBpxJDbgPoI+iWUedjwJ
ki6mNmm8rrqArDl1T3lSTec14gslSHooAlgblIqc694sB8jRcXlNHFGenepnBvSEnYw/Ebe+XfaQ
OPY9C1xVS8SOXRXF+yQCVWxXBsLE7ue5brEfocZQtAVvqEcWqVlOGrYT9zXj1yIzqHkbdtylhmNO
ycms26MnFZEIdB2HbI2VoV7sysxWdoQ6qKPoPLD1j3Ih/d+3kR1TRm7uySuN/Ld3OnMx+l1JjYXx
89yYy1uk2PL3fAcBYpVv13QGl+h3iIYJBQLqBRBPID8lYZdAoom3H3BrRf9aPXSmorcKp5iTcudx
7dBxzRyua9/xLWJDboXFhTUsaKx+zL4MT663WApwYQYiQCLbEn/C33sMLTiZVhKxooRU1peLD2cW
6EYLx2UZhMb7pSuWU1kZAqXXq76b3gsWLq4fuu0Cq4m2TFl5wJEWAnaLqYCyDwXkCiuAWqgvhuOO
KW1Xr/iWPutrPhkCeQOwDcMJvXuWvgzO+vIB5PhbCcXjtKkRR1Mf8g8NwK3sU2oCOy1S75BkSkG1
UkI2ZPBkfzoHyycugZCltAnRysAWcjsniO7jdWZnIwan5xEnO57TdXXrHXYkJn+vma2KOzY2AA8g
v6fhw2sb4FvDhveQexHeOEd6STQLf5XgOfrHqf2gNfzOYGuVmNzOc8pBzEpMPJxyTSVzFeiYz8Gk
ViRakyLpzxLLhkn6TzVzDPiDOikqfHkUHyLb64cyEZue6TrZkHdyn7A+HoV4zvTVPUAXvdF+WXZg
mGxaNGA9Uz+YxkjwF/KC+jXWP2tHd0KJYVK0AymXBlSAReQK4hsmUv1soqR6q/fRaDG1y/9N6Z0P
VvGHjzYKOGci2BbjM9Dr4EnoNEKn9bdntIUyCaTRJDUk/6C10wM0xtSsWw4qjA1Y6hNs+zClsZsG
OnYqghqVCzEZUKZLigv+9/YfEvw5nvecqb/07LThdUalHk3V+96Gk7uQNqJjUhxS9KATXD3HVEt/
J7GJ58tEv0CmwuCcA9L8N8c4ZVWk+7GmQ8hQh+KYPx6XTaV6YKVrUF4/jxxVmT3tOZIO2vKymhKy
VF/UyHd8s0f/pQyYV5h+eqYu+p4QVFp5gygxwh5EAnOf1yQEMJyM87jbAuneR4v33imucJeBmVr/
XMTMcmvpX0dPCqsv5PcgJ6ux6rnNfGGk18VifV6cK9TYfY7V7kd6ctGVPWzN9N8BxUJUdVgXcCOG
ciBBwEQlwnFZW3DuRxoOLYfsbjl7Numiergq7g5cbFvD2xtyohyenJkrVVVwNhLK9PZ4AZM4OgVO
jBH4ColTbj5+/qdj2hwVbghgIMhwRDewxL0sG5XqiHk0lR9SSl6cEI2XS1iU1wjaZh+xDl7xfpjc
Gv7g5Cz6tisfs9rLPBFapx7IYtKVtg4HEUd2jAuJCVtP+tjHcdfqaKfZrSNeU/dInMAuBUKs9U4H
Q9wYWvNVn1FTfx5kAv4RlH3gV3dgdkKRw+dtVsoiBRudd47cOPM8z0m4BpzQX9KJxJHdWHVJByLr
1mhoVttD1jYJ7BwDPQmYXE13gomT5PrmuCTVfpZKpFxU9b4KszBP9TDinPmVKcHQN+AEM7DYkYUQ
U508GlD5qi5oUMObFUWI5yb7pGzkw0EhqiVPShu+WhhZ7ZXCFLn5WPc76q0Kq7UuABDcmrjhpkVe
5aRTMniIWkZsEd2lHW1pqz4+tihLCh7d0wcHG2JoZ9crQge3uM60ZeEoZt+AGJjggo4RuYYCnJyJ
O4fUcZZrXE6p/0BKRK8I3lnFOoMcMjZTDyZsEyMIsnjjGBXDdnNY/S8arT2xhy1OZsK/OA4djqSH
IfVx+hDOAh03S5dZ0zWgAkrLytUM+bDEfFOkgYX3YwSZndVO1weRvAj0iZYiHqW6IHnyMAkc3Yrq
aM8S3LgJ11x1z6ledEc+1074EjWZX7ozpZsjXHWdrjkBlg5Yqu9uaw8Z6D18C74v8OBPU4llj148
ZkiPVqusGp0CmaUpkMTtLd4acEQpwpRdjbpAgjGg2w/tISCFrtnv2v472yYyhbSAH5HFkKNt50ic
0UDhUX6o5Li3Tr0+WPDa+I0LZziRdpWtKatG2qkB/4vNHfxesx0Wz2uTtabUz6vSnzpylEFXgl+D
WKihDeLGqZt3O+nUKTYm4mS/tS+AX2sZERfHdAqLhAN74MB+FcKRvnCQpSJfxMCazLC6ASBKqzmC
4knqE5sCBbusBU0eWePR5JC0Bf2RfuFSn2dRrasiqitAY9S8v2PdsBX34Z57S+mke5vA7BbglPJi
7P1PkmAjSZI+QUR2TqxjXiwIVkKuYh8oh5SazqOJ1gUTCVx+EQFIQeBaaFjp/lC1/z7aoBgzjsLb
0Jk48nUFQdalnTH4dwohvVvGQXH8vvqEVhlqeYHmLXNlCTtXKmFJrht82DJTLUAzf+275e9m5+/t
488BiBbB2A4GCDdoDD17TvZ0B7aYKoQwcADhVHfDEst83ArUIbP9c11r2mGH1vbABxbHUJu8aQQ1
0oHgmRD1SPhm7WYZ69z/NUmsVNwaKP9SBtg0YwOVYggBpgkDAHXVJjvxqTZeeLiK8SV80mHHnnzl
EWgMx3wFUVQ0svx8/KHUXqR8fVxFjCz6yID9N6Y5fzdZU/vy9Zyqahf3Ke2xNBaIHbzM7o1zdbjl
5xcBrRj5J3f2zwgEluSFILoCbSct4QcnIX6u0HdE/t2AdE5Kvxznu8ltxHVbAX4SF1+HW6FAzkBF
8oWWA14yBlqPooS/XXqgKIX02TF5VykBq1EUutIFyjUA3mp9SqZB1u6UM+YRe572H6vnfLJcfsJM
H/wP0NdqWPzOEn3SuK7Kqf48qBjfnTFeEgx1G+RPpDLQpH3JF3TlENSHZ9Psypxv7XjhP4cW9OCw
zYbL2isgY6VUyy0zrObORoZ5ovFwsGA8YRNX6eWa1/SzSgOD1pzxfBny+Td+vE3CZqArXe7EKuVJ
vinnzeQ2Wjw5NdHTeE4mCZj1dA4T1tlg8pm9SVsfF4tGveGvyxSsJAI7B85InabxhG204hIJcfK1
8frzHBxWlkcDZdwFvcnEhAMmUgGnLcTQS3+s+82bGCYVnSvkRHFLzoudcTw5AJEswUXhUQvht39g
s6xTnuh9NnuCh9mr/uVl0yf7XP3m+p6KoNkZdvjrRqs2mynwScNSHUcbyMxC8kPhyG5nHdhn7HXM
Rht4KIijTKD62ohfP3+ZTEtq/D0q1roz8h/gGYwefDu/1bVDAa0F5iH64Im/kb0hoN+l0h5GSfFL
h5FtX7xaUDZoR0E8HO9kBg+T5l5qBbS+m4iABPqNFPZR9rE/0zuCCpo+pPqRJNHCtN1K3YRxIDlS
7m0AeF+G11L8rgCRRtOqeE0B1bP41+JbqRowKsWcggcMtPBL72vD8Z/n9D0UT9k2E2/uIw+yPd85
xB69aEDPjmUL6Vp9kjCVxUk0zCk+qwpj5PNaNIgifpD4aJYUaXaBq9ZOiOTNNFwN94TG7H9ofZNq
Git7QzRCWwvjzkaB8VRbhBxbUDzWX6EN3fb6OIYd6Sw8PK4Eu5zq0uJqPiYTzFrs8uO56FiHbXy5
saIFn7NzDBk6cKLsOqGxjnOGXK2vWqbYbHx3C3GiHG3NRpuy2ez+L2jfkAK0p6I9jUuo7JH02Azl
B2bDSK04TD3+dPu6tDR43eO1WwPCCcqVEnouoDsiu6SktGkLjxytVO4Nawr+q8vAc9nxDQBXt2Bc
M6GRLYttjUXgYXnc/Ap0wFrBq1eDMgWTjyKDsyX7dVhyJc3jUiHeirvAJN75Amg0rso3FEGl26vC
/gTMWoOkZ/dGawkayQljcla2//1JLDYOXeVCvnFlW2FvFtVdU1VSpZA740z4s/+kSNWXYq1lzuE9
YzHXRBI3L7tiewEoNuwXl2WojLOLEYxXwB0mDsgf8M4LbO04q+4gYAtChWVcYb01KGcl0wn2+XFA
7yVshq/zNbY7ztdUC3u2x35634pAk0193DaMgm1EVB8+b3MNiOw1os8vQT+1ehquIlJ1bpmwc77U
Fu+tnyv7sJqy7dcAqP/mcHotxlA1rAlo9HLkpJ9flverYP1ik6MevpjYJ3Kql1Zs9f9deR0x1/2e
MbtDngDqvemeNIShElgwqCzC6EdzVPIukQFgy4VPeDBBLv4neFwxc5SHZpB4nxS8KDenjd3wAGPl
Jrjs3HcXyqm+TPp4NJHg+VOz6fDReHCjKdsp0OocHkTENtufcdb51JIz28CyOu4DijzmXAVt/a6G
4XNIzNUbe8M5tSItKBWy4asvtZIpUma+pShsWIuk4WzlDAJ9zmxtYtSEN2jgpkDzJVuVZdrvOYoR
jOqOflJXwz4JZWPUOmC1XaK+mApBp63KXLXc3ShHYPBKehqz2PvTFGeXr/unAYftHgRdBmAVz09M
P77koDrQ4slpLBTwpQbW55u2BaSmVFgOoXlAEhwR4WD1yVX0sw9ffj9MXzhw+I/ctMVv3Dbvks2R
Ke6gOtqp/vvKaXiVBk2tJh0nrDDY7bgaQEgmio0VlpQfxW9mUPfe84jzlxqeBiCsyK9acVODnzPa
iZ+dtuT+X6k9JUMQtalkhiCFzemM47RIxRgAdJYmQU+i62uLDp6k88B7C4Zyu72H4/MFDVju0oi/
AqOVJliyiOwkX+BtDsDtpkxwvI7X8hhn6T+Iiw4IKo4pkTVCnEo1WL/GgvlfSw2dOfbRBfYPADb+
FQywm7dgj3Au65xiN1e3My04BSGlViMNMpqbfntpA6oCl0oAPXylgAUKgs5OeuOCE1XottIHEcQG
6waaj36zfctoolKbgxOF2RTCZ1GDY/2p8PCQpO2NdIFpnKef5UTvycRaDebSenb4MdWZpwwiWHAL
+s6QAzs2l3eBlMvU+tgYATTFqebIJmq/Hj6aTlYnT9QBgBXY4rl7bJzLcTZLZ1e1eR3aZg2xQQG3
RBKOIbtJsrx+bUhkGxDJKvnL514VK4mWWo5lop2+PwSTP2jZ++rUy7NSMt3On1igbMHZahbn4fiS
2AUjLxaKAgOgh/PqOa56DiBn7Sr0IWz+k7Wqsuz+Yi4BB90JtbuKwVk11ZsoOFU5U3esjuDsi4nZ
eEpA/NabZgR0I91Ythhvw7N6LnXZyRIJWNIwUBxXH/ER6JM3UUtAcFEAk3PwuaQjZMAlUwK0LiVh
957oDp1aP9TPDBd/5xGqNTZbSykgCprxwUWB0TCibSFRUQUL7ajuHZc2kq3xXVrkUp3/tFDJGMEA
aNIKVuh/CqvK0rGVSdYGPupMyUImfqeh9fjPVMwrjlkuC+EtG6AXtshHBmkL29BDV3cZbstMS2zt
S4N+d83z4RJHrNJTIEMu/qaZD/3yJ6gY7s7MtwSdpmiioopo3SSZ5GESNCnVbZYIp2GDxpiUt8F+
b+FSbvvThkCbhGtmNCpa2K/FqPTccYajMXeKc+prSNYxejvhtMhGCuKguinuEwO+KlXPPsC5W5cF
zrFsWmh44Xm1Za/bYmP+xBXJz65zEOkhCMoAtFKBPGGG+LK7gscifdC0a0P/u5Wa92sfRkZFl9/W
YTX+CR24cn3ezARwgwywl+bw5gbpF4c4rFFERM5towfaSD65v36znC2u1iqCfxVwuEt7fUZpyOPJ
TZmVDmffeAU8zqI6tMtq94uF8yhpoukSdFa93xLNoCiTWZsgKtx8/FjBEYumT24z6xL2pGKIVQAb
nucmOOJstT3WiHKMNJIVb/+PaoXhGWEV6LEu0jY3eVLYVHMcTlXHXIgKFLmjXlDiDKQVvD0enfqE
dZQPdvYnt9ChGfmd/yJfb2hrGgnBSZvzgQriPMuxnldoYtavmOHA+UOT+WLMvwevm0jN4XsE2+QD
d289pU6Y2VlosOFDUuOY6d/OsrncDmhQ8RTVfAtKzsoo9kBSz2s7VShnWt+NfcwnAuYpo4BzOoj3
8ReJtMfPQzmd+Q13+wzk1isB1ynXrmtV+xKNNeBC83iwdCbZuJ1DmKLLOP1MiJd1cmULhs1qyiuk
yDHSvVAInv6NkbBS5U9yzO/wVl00mQF7vhRvDsE8q4NDWYGHS61uTkApBSZZ9taK6bDgy7ObjLOI
+mQV4UxYOr2mWB/5cDv1lBkC0+w5RtzWzWTVeYZzMHnffkHBVqYoNTC9kUZMDmK5S+u7LtdhaO/Z
ERPtrIiKZOGlWL8Jk7BlLnVxf2L6pMgiGXW83D7iu4C/yx7nqX7B8p9OHCagGnhxH7Wdwu23DQm7
wwZ8g0SsTSqDNC3FAUKffmJc6MUl04zW/ZQW6tuInNqO3h9yvKfYBQiZay8o3JiD3cc7hRbSdAOd
Bx6yUmV+JrqLIkgdHEHLTD/Hfoiti0joYrCwaye9NzGa+nkpwWjjNYxqwEcEkEpAruFMVl0SXBRa
RQAe4yL0diybrQEAgnKkkNMN5p9/JPRFgNXvZtVTlSTLKnte30CsTop7sAcvFd2wW60TWLojdFt/
9qw8u+54O1nK0PgcC7Hdl4/goRoBykxNGjLfwBTD8ut2auPnWJaYBoHxWTFGIOOe3SFsdgFS2/1D
fEFNm8ecTp2lRQq7OG3Oq161D8qMH3GxRp0XulXhGYZEq1a6/EJG2ORflpkL7hlW2Q3GzeRjI5r9
JeoOdW6KZBqmYHbwccA3u+q7JYSyA6NcuD7obQ+Qcto1hN64fnS9rc9Sw/dHc99Glf8keKmPdWrr
CUmyFzfkwDZng8W/LZdq9x4w3t8ufvlXazj5axUoxu3iUNxe2v8BVTzgv0Oo6HdQPq632Ep6FGA3
oY3tBRC0EMDbvCCWRXPw+LQFzZEriKrS92+h9gPEzg+XdabSlTHUqVoyflXLdQ8i7/XZHe+iEk2U
JnrZJ080hVwv3vWUm6pK3EZdws9AHrBGYTc2z9Quu2b9axMikOpQ6ksMQKwRGCxKRDgko3LCHVkD
Ko2sRnC4FjkSCZlYs3TUooVWyuemmWvo3pmgJ04K7WMVkXoawDhIrFJP/WoKEFavv0Px/CWYOMzW
KhLue3eVPuXP1+BFtrq0iurx4C5HmPWeHY/O33uT0cewJuQOibvubo3KZFmTm/KZ4h/zucZo1UuG
h1JiGYDZ3FEwVe173zpbugbl8a1rOvzCYfRjaq6E0Vi3z+O8CnaIrSeC/k17aVQ0mgtR5lrLpLdR
2EvvIoZnJn5X8fwjES9EBGYU3lm2Aby0UxT47V2UlreQc8p49KHbFWDnOeRjMuT8ZKIrYfdcmWiM
4LT+H6wK0d0ow2gfRmCBYlI+gqsUpgq30GvpZUtD+H3Z2Uuko9rCd/mBxk0q03YYZcEeumoD8an5
mBkp2DqrqCh3YFrHPI+bciQntt63lTEn4BZrvrWNCaa7q/9rRXU+rAH0jEi3yD4ko8LSeLCIR+Jd
uhdn/uYMavs1tm06J0z0KzjZawplZodutG5JTSkv/aykglUjihxFWGbuk2k4lMIyup+W81egvw/h
KFx8AKGLBJd5IaoeMJU0Iv0RWaxjK1q5J44XlJkk1l+RrryD9idtMTBN3/sUf+PstVRWKHE9Wzpb
G1ATz0XAiUsDHYw8I3gcfQ4wCq42PlkoQkZ+9Hh2NRD8uMNYbL45d8HTBnoWirRnuOaPj8/0QyHz
w7iX5r4mUkIoCaYSk9t75XVM/tzzZftzDCy5apgU/4pgzwssxw94kTHF5GmAXo8SvVlm0a+ssQUy
8RYhzeoMqeWKPiSf5AKLImdZ9UnM+RG43B3VTfUZAdsEq0D3HiBc+pfk8PKqjk883oE7nEcHO3Ah
3cCWnM7s9JMPS7tC6ZU2fVXekdS1PaWxQ7w6Z3thORDE5sy8HWMoGA8ww8KBt/kpkF04aXasx9kH
fKaVfapOTv2iEGWrqq5TJvcm/kgfDgLRpWIclMdN8TG3JmqAITgUOvi9Ht/xugS9yo+C971HLjwo
WTo5C2XnTJvPuG6cK27f0obJq4STLShfNmA8lnmNeGlYnBrmTkfl8b8Oc17JWKRNbG/n7VdPA3KV
39g+xoYoyR8whpqgJLvjzRQf2kjCjmA4ijp9khkAwk/M6fI74T3NcVkyCUSzOBQnvL5ZsPRmlvJ+
vvBtS1cgl1+e7geg5mXhYE2QmaOn/5YHA+STXESI0PNf2lJyCg3Ot+Z7DWXizkq4QIrdwBHDL1mD
eodKci94PsECQh9gx4pIQ2spt0Lu/QNchfI9xOFCX8+S+T7QYZLYUaRPuNcPtoFgKHlaekTRLqSg
a8932hRhiebmaUgcSkl7ZDJEbF7DYzkrOOlgwt+dx/pgNHL6iE6lvsUFA2Df8ydg//fYtHNez8aG
OAYU+Ls8MjlTUi3Ns54MfElKeW38/YTO7AiQg39CIdQ8xuaeDTO9FJLhgBzVOZuUw/G6ol4ICxv8
ZJel1EucQ/o/FFskyHoqLsTyQIJ8lWVATuxaajOA9o1TR46T7fwp1FmgBIKCj55sCrDieAR1uuUa
nQlBdEYYS1g3gqsgpq4DemR7SIhdSn/K0OjM2bsMKlX9w93b8FimlnlBtQv0Fp518zqWw33l2Rmd
7G+ZHIzp2HLUxhe8dO4+ibKutnynOoW395DsgrsaNwz3RrJRoetmhOzXGVFckoSQD9HaTZuiZ63m
vBgSY+iCqW99gTpYx6OfcZatZBekANpdwtap1FAUUxgWmn+gb6nINM8EGqv5vRD6jl/aBLsZ8e+n
H7AtxpPEGUF884YQqbv5rtqXIRxjHIcs1uI4wtmr3U3wB2rGt0oqxE97guKGvYzhz+PkfQN0NEgK
W6daC5aF076E27Yxlqz6LWaiGRpdu3kT5QmyeJrtH/mC7MDBOnEUhAs59ZkuzbTzIiRoqYsuK8xd
FbsV9cOi95bPMg1CkcJrdESBgXOuRjPlrFKd5cc7ul4JhqLcJGHtNECaGoo31s0Ik69uQFDp0jmX
HFlGr5ldo5KuIjLJbK1fKH525VnfTtQ5GdQXQ+TiJRL/SKmTq5Y5bAFZCd+pqRn+3VSjte/UTqZ/
gMR664DXvry7gENyw1QLxtRTt+yR3s1binOPvmIcn05j6SC1kHKB0Or8a+AXqZPeB0N1lMZBBtl4
8t7isbw2zVgLk3rXGsQcLQwl5DjqJkcbl4BJLI6bDES+vTVGS1QCELsjr+OCmgJpDmc86+TCQzkA
AlMktkI5oNOqW0WHe3Ig7FOWdbO20kOEc8kV+Kkj9UVshLR3gO0CoeAH/sxe16MfFrncXof9Os6A
2rBKZYurhrYFs1izbmrBQZdUGqzD93W2A3cbrvIkTZetgXSNJP5Gk+DA7BQWpofoToiQQJZApY2S
fX2/ScWytASLeBjiIBkfH3HrmytSvJjVV/NlfApIOdIyHDsfk4Xowoa+WTKeS4rucx+Jv2l4trDJ
gyhTkb1zCQYbl/Rsnjp+VUP1cgEPOGj/Grg/xqYvWKDwvuvvFlsapl/14PZSw6/i1Mmb5DbxrZYS
BvJVwYmoS544afDPBzlc5r2Qx/htS0LNeae6XHzbZMrEo5mcp6j5feQhPeQvzQncUoszhDx/TJMJ
fhMEtT30AwdxS9JUo50Z9vT7yDEok2q2B7Sj89Y29O1q9tejUaLT9cu4kgZKL2AaS8hI4WxcB74Z
Gz9bLYxxThSJZp6J7qtys4Njm8L8phofgrtPtqBDihl8oPqDQCiHMRaEMt+ZjAzc6b7GbTBEeFFn
S6p6gxBpVYoOhkkH2ItzUE80fgxW/XwEva37a4d7LV7ptv9f9/HIhoCNyiHdnZWOs2hH4ZRABZMk
6IO9hFuOmvcwBpeZ9i7Eg9F5RpAbtMfwTdNmdJD/rpklEJQXKgiFJBlwYLyjHdgqmG6q9craCnNf
56gai7ml3aS3qdxgQz80ZHVG8dE7Ipzw59GP6MFC/EPPVUanAzuD1wRJ9uMKzrlTfLJI6Q0jDZsB
H6V4DUC1HpXMzJp6Jo8rxts/7AYKXSKOvvJi5RJsn4rvCvpoHsxLZtbJpHkV2a8apngI4cSX7Wb4
vGrYj7PlGaWAhgR4nPBPzl4Wl5MvWD4OW3pW50KH8gh/zOerV9yONX4NDYRnaZofa2d1gmo4DnFD
L9XEuxIB4Gv3roCCF/wQQFX1ufO0QH76vmH4jmHA5niB5qjRKFvk+wcjjkRFwimk0P9uc7icjWlg
yzoKQFDUjRX0oPeV7Z60SP8uxNmGn6gWRd2Rw1vyVIgw0hLRgXWloE2p4HZ0j9yzSySN6aof3uRw
76b4M9Zc27wg+rV18HciMqhcL5jjZKn1PhvxSzK3nQu7B5rIEuLDHkWgUiyqtAjW30X+dUamBdao
sjx/mlDXIKYJxtOeP6/JzLXymG3oFM0Y6Ihy9ac4XUJXDAS5pt7CEhbNq5x6PvN6vDuOi8NXjqoB
CeV+95OAaPePTQNOAPu951gmUv94kjb/hU3RHtWUE7R2N8k9hVzHb0c0xoCFAhlQ9T6N0Hhft4Ks
/d6vKkctcBGAG51HDyr5LIrQ4NR4ZRVmSxb2LksX/ULrrZZPUqdsCBRIEqgRfmpaKE0yfSq7+WIQ
gIEBQMHz/wKAWtQeuMUWfsF4tYpVOHgkWTeffFA1YhoDkEwarzhfkcSlEidd8J7JWwEM1FKX9N7M
cFgX89AvFQdIa1ElkIw+jD1YW0UW2j3rRn9p+UuPplWpzvByxf02fhWySImrAWZFuxOQ3TAOOZG6
WfamEBQArGjgxIN+uq5teefceQ7OQ8XZ2LfQieapaMBPpV5cb21LDGR7kV3fngJMY8G2tT9QMsB7
nnIcL9iorSKuHe21XRIx19jpTO5HUwTf58ELXuvkIaKv8myhJl3JmD9qzjCU8Jk/xcZ2MZfv6xWY
NW4KULofjecFZ5T3HO2FtzxMVmOJ7MNHi9aJtvRgkZsf3KUGbE39b4vggL8F3CW/h1KPun3xR10w
cUzaBMjH44C2AQXxncXOZZEeWeHBsratKYCv1qbOpm5U/deWja74xumR0HHrvB0OvMKxYbzsNQd6
ZXzDadu9r6TT4TIgAlRDSqSZxweiUVuDZHMPY13CsDoc4Oj8Td3KFUd9mw4k4J8ZkWegbbBgK6g9
K4KbqKPSY7Ohi2ui4ZxasBvrimu/0MRJkHM6VMVXtnQraUVirSgCEUz8A+BtUElf6wbJ8xnd58T0
Wljz6ZSV5kU6WTP6/yjnns2Mge9OrBA0RXw6aMhzFJfod/zY+xafXpzuDx84dIvvPAbfGhz8zlUz
mI4WVO0hz7EWFmgSN3cb1vBA4kE0QQZYOtaE9kfxk65gfUBgCSbw0XF0SwZuUZ3Vi+6R6ZNsl6+a
Op1zZVtgjrhzlS7zo1xk/1xGUON5vgK6wS0AQNrcQYKVJq1a76+w6/bi5b+G8b9Q9Kgel6idRi3+
5htvAJ5EjzepnUj8ueMTdhhm2BVKGt6IGGl744EEdYtu6wsWrRivaVf3OGH4rpbwZeMRW/PgxI7j
1lmUd1T9vkVl/4JeCZL1gTnMM7K1BCvbgai7QJfwfblTSMZ1QW02nQclWm4CWCM/LUI7Yh0mzABl
u7T0zJdhC2DSiTU2u/pMkYhk8Vk5obQ8botI3y8+YvzEEKd9HajZGJ8KOUsseWkMOlcjkOw/6oJ8
D5Vzms7HCeOS56l3N0/UrXvn5mFI2+hGeF898eadcncFDZP2A8knUV/rI+QFFfoAx22YH1bTus5S
kkxoODZM1hk4EtuGyO8cPkgu/Jni3jpPIr3KyQkapmmOqk0vfr6mcVkCJiMvbvgEbviHKWXtJOZg
MWb8YKheUfOa70aIF1qAYZcoVMuobGFpG2cJ5yL+n97hKjjtSR415xJpQYq2vYK9BDq5WJ+TQLu1
kDuvajyGUsJ1fMLp9d6hxwQefrp9f3aKeMGXDgKQnXIqXg6n/BwkcVR2v8HD9i6HF8zqxSjbc9M5
fmFqRaB7fcI6oXpuqT2pBe8TvcU45k/Qk+31Yk6bBUcSnGnPwV2oZOi6KKLVC3ddRLTRIiMOeWON
CdDa5ePSnl03NjoI549cvJWJ7cVQlxe8zA+qwk8UjjC0XZ4SfhzxVgMSxMoHEfzwoZAYOHjLYUHJ
sBq4kqUhF5+WSD8uijs/ivKyrRL3pBShwAt7gY1GtbAYCvvYj+Eh8HVrmUeNei3+v3/fElZCj63J
WegSgyKCnc88vsVLGPa1r9XE88GXE/hCS1X6VaZ8NZdThlbXvXTBAZ55V53WGnZMTVhKGxlk8leG
zEHyef/uxCaHMSbiZFcYCZD2uAEI8Axa9AGIhu2y0SSuCFWJd3hlRFtYsTCxPGZKudgMCDgTJusW
3zm4HFaT1CVnkpJ1xxzeyBG+zHuFHlOEBthmg0IWgxrwaaRjISzgEcfDYMhCcgljQBGAyUoAq2od
EZy3ypt63W0nhcGsb12zmDJB81MpbpenM3A76Lj3kHZr6+hXkkkna1izBrfcab2c4SxUBVTan4v+
NYuT72bxU3yo9sFCpOln4JjKSjs8RhRkQMS5WlDxQwNrOFEN/K0k+6HcjVb1EZre6HtQD+5DfNFv
h0sxxZCiSMyUUHvOjigbQAcVuGu7YdG0lSl7aAi5idw0kxC3yCAvubTNvJtZXksSQy8k23qYBHY8
YasXGTwRMPgfU+tJqbM+G9hc3bROqNLaLFefC9iN8NDaqCdB3udf7s70JDEEGhN126eiHyGJX0SJ
PtT/QBHqTScYsFhXvx9gJeB13Cxv8EhiuZevA6l3EpDp4CfsX6292J88UkvpZ8kt+1C937kAASZe
xO4UZK+ERIXkAarV1+uqTH8QOa93m07KAJZDvrL5JH5Ttv5otgH7/8z5jT7X4b4974wthvI0zlnL
bZlpyDOigonGmBwe1Sbdu2O8kZkzYQ6mKkEkqQR9Qn+/tQC7zyXs4t5NoipO7nKU58C8xrKnBo2A
vvW4IIOpqfW49ziWh1VjnMcUA6lUnkrCyWcZyy+hHcihct9m1gyb92ysOUGWfqYWOY0XpAv8TgNa
hN6JyVy+Kv1IEFvrgenMDUeQnJ4zcvVcLtKn8Jz752uy3KB2pLq40NbqI1LvN3XtLpyaBDlSdA/Z
jAOPBZFvyUNajcGLAmn9CJg7mTNM1TnEpWRP+8izWsbOX1RZhqjgGiDs4YEJDzJWF+s8hxU5jIN8
XHWXK4dYbrvbVK2+ce0PrqpY/SGBKIeCORBnxEPgX+oFh3ijrQgzzIGqmoRZpcNp6t+bN9MAOl0u
XWOrrRTEj1C7tZT+qsvL59eaG4tbz2scMr98od/ooP2zLCvyehz9r63OXTkQyo5yzky5BUtqF8r1
kpRhO/Oqj7mgxd6MwWqD0aYHlhlFGglMeqe2kX2x4gDpvvKXjG1uqIgP3D7iO9XtbV3QQh8GXnHQ
ZVNHF9/x+F3nRP/n8qoIu3ioCSr8KE1xQNLLC9k9s1b3maR0M22ziZqLttneHbQn9TUY0j2y5xZz
eTCRHE4Vhfvf9IhSAPLlKzfSkeOmZWIu7HfjKX4iEVxmfUk3bOufImEDfhvMTrqJ0B+9EYf/quxy
Gnd8PtYvQiiA0DfdWPjYkgB4XbuGZu5fsdzESnGe7PcMm0yFklshMgIUNd/MLuo2XSxm10PC9KsA
sxwsUjrj3pV2WZyw3vsB3C9fNxfL5/laCQAcF18u4rJTI+RFvB5HE/FwfrvtLep05VJPuFLLuyZQ
w8+ocSz2UJgjcebIfBxHJ6ckATQyrbxqSL0K5kXk18sNEUDuhCOWJqCNgwvL+9PccliHociNJfzy
vpphB+RECZhZEy73KHVyGNqYLPnI5xQZZIeZ4aBEZEhi/mhclOSIuKVnvD0LMynNlXCFX6phjghR
XkDtmHC1qh6yoxcXszpX12SsdhQ7+iYrTeDkrsCaqST2EzbrJ4+Q0OV4JDsiHRC7Pg7BdvKB4+TB
LT+3IUCznfVNlcdFIaPUSmfe2cQcIfrAfvFttogUypvKfVjli8TYD193HJKxxipgUJjIjozC3mom
m4SACuEgRsbrZN3UykM5WIDSpQ3/rHSiuXzUHBfzRofXwH4NoFpZBefp7Xrj3F2vGlVbfEelzh0j
WhwuCMlfbEaFG9s4miSSqZBRTNSc0RoE9Z7eGHRd35JtYXQy0H6QvbB2rHROLB+iJjGqp720MC+S
/akOcERSvTtA7E4Ucp1BuljONdd+uArYQbhwj6kWhEXnGDTa9oWN9siuUgUit9AjV5Gep5IpqC1n
2s3+5QCGpwfasw2DZkSw7hRTAUlnVA8iBtwDJysOoYBC9OQ3VXvU1o6igyOhLmfITCcwKMm4k+cl
KJ4pfUiuLKrqFw9Hy8mNFXxJ98XKcE3cSLszO1YsTkFqZjxjPdgg70S2wT0BJRUzAQ4HNgVZftJr
U1GOwXlYP/LTnoPtW8NSjSvoawZAePfFbKGZK3BXrfRfywY8uJ4UWcF+mN5FDUPW6qmpYPyG78GB
qwNRDk14G71WaaB/2M2q9Y6Izv3Y3okcpE8y5Pmj2Le1ySlEixlghSr02qurDh6YKJMrUVBDvwtE
vpGG0XQo81emLomNfTE8I1j9MfLt6alcncqPoblYy9/zzUOsQvsWBRG6HbHbAhbA5PJJ+uznOlpQ
0FRrIFp5ezw4iytZbLCh6eZ+fPvRb8TDwMWlOGlTFtDC6VxS/mL6eZZ3PtFFEuZpR2IOK/4YAkbI
lQ1f7KPRjmtbeZKh1FC4qNdO218NNaaASZ0+t0Ursel3+VB09VoSqwSrFzwrE5SNp0aMJmXHwuTK
ZNpVivt34c8Bwz0xKdRfDT9Q/irpbCfVlYl5VQXK/9yqbEzrTNA2346c3OePlRgpxwiPNWYrl1Qk
rLv3MSbjWGD7lsg6cxso4PhK+xuxSM1Q63Jxb/3LQflvW/0UBvnOLoPOctjZ76Ywtjwzu7shJ2BN
jNB6W2P/DjAx3S3WzCAKywEdtl95UQavXt47QqXIP+i4h9FKoV0YDLHdO/7GhJGf/NkacZPBGx+/
gmqsSFor3aLHnjcg0c/xue0BFiWsI8LZzC11iznxQhZ40hqiy6aHu/UW2hs4NRffY4URBGgK9G+j
LfHb1Ck5mOq5JdfYdkqlE9QktLp9dYQ0uQG06vYooYzAztFMgwGBW+Zsy/CY4leqJNo3K/cfKI4T
fZzY/8fvkhUmCP6f7cKyssosyA3yLsFxzSYym6LMcC5oG7G1JJ5jCMHorhAXEB6zKpF92FKGrs9Y
pMAR5llDBFrZOS+Ry/I60ebaAY5MK5obc5i96uHg+b/LKL4YOXBAgFOuhrlpdwdeqOrrysOtXi6J
W0K4njRcAKMwbtOCu1GyW4/sRGHRU+KyVG/hRQ76cia5LU8JsbCuQ3eSAEfGd2BoFpXAP/hfqvHm
dAb51ohkwSrmGq3KKSR4QuTRwVMR63eiIgBbggFsFArnCS0qU4euT7F/EzoC61h427ojkD2iyObS
4V1hUgbdyNbyDspECUwrVrpuNo7eQOuGYA46tfNX2MduBAggr9F0Zm8hUVKqxtNtnL2afovwga2R
+AH7oeVlQrT08srYvGtLwwX15AuTz7N7ft79h/yohGsNiB2SSyP9nuw3IjYov8eIIzcj8NLPvhLG
inhC8NgxsvDsQ87BRs8RkMtER8+TGibilm26mReKOXbSOpHz98LkVbrmxjKUYcuMjWeS28QmWIQM
CbYCzxEJ7Li9/tmDk5K/rph953cEwTxMULFvXzqBf9IouV04ZZxrT0QdoPN3UfSbOSFDZFCw9Ucg
NDDRRYsHBz90n0aRP/EdqiWSOggouWjOXctdc0JrsPqqUp0jQFI3RjYLwk5MzsQi3tu+t1BO4TbO
jHzw0a3o/eGyme1URDSabwhTiE15h2yELGyQ8P0etyoQIUf5GkgY3evXifxEa0TJ533yoF2AYWLi
27EKkxtnLu4j9rQnAxS1c3J45vFU4up0Vw2zovDfSz/mRjdwYIP+eV64q8pNd3Xd7eCc4JBaGCii
Kun9Sll0FtwuWH9As7iZCLGSI/54z9o906L8UkPTsCGhuHGIUfxx6Jzmznq0BXYAXtzeAzZmr1Vm
Rxb3bnzsZp4qMN9EoPKE4On0HKJeu6r2sf5IPMJf+AJFozUbrb6LDecKEY0vO0ziAJxooyTIZDk3
5w0CS0AlmV3KOECn5/DQQg9qO0UGMXyxbionJxMQuqraJpS/SfexHH0gDpzRZr1eb/IDNtMKHPHo
45cEPF0GI0EpxrYqNlzHH2y5Aj3pmRWSZcOH8j7egRuViCLPz3LJS6qQvTV/G68gABZD82yqdWPH
cLb8qGzbxc/ajcdwnZRbzLEts6jtOyksTH1tqBahv8+WLJTB4OiuLa5Q6CTkbeyEaGZcwXygMkO9
MRaiu8gYxMuAV9CTQpPm8zWhlJxTW5oJnHiskxggxdOjifMbN0UGpUxD9vX3qknAaxIpCOjjzZ4o
OtTCz23n8E4sHY1w6bpslGt/C+7cio8PVv4fh7VW6katrLPg06BoJa6wnvklJYFlzr1gmRaOGKv9
2Ez/iKTiqMQ0w1gmQfH3Lw2OYfEATPT0oWxJL9xHajFaLTC+tD+zdl/u1wf4pU4+QM+7aj4Yn+Nu
Zsri9mQbyOjRATBHhAlW3iSS0Om4IsuhtxPv5D2cJt/xv4A2NTnxCLQlf9kqB7qhrBmAv8m7stTB
vNiJdgyrn8lzfkKzYtpgoYZ7NAqMjsU0W59+v4JqvE0gzzkDBgnDtGxVCWgaApAF55aGUND43NXy
2gPBIT9SJ1cDORDMzf0rYy4C/2Jb2s17asOl24z8ZIkZTJJBPAl2b5qldr755h81LkHiW1BghYLf
UuW/QhM2MvPzHKuk2HsmaoXEPhULTiYIFNlb8sl9uqjNByiw4DC8YTMsaG24yefo9dsGmbOouphw
TtFFzWNGW0ot4W9vtzXpo4g0KmevS+PxffL4LqcXL703XF6KpAv+tMAsyVB19ch6MPEaKMK/D087
d6IJesi9BgvaVVS4Wshnj7UPWLRL3cfU25MJ4HfZe+hHpYnmvIrX2xjgpw7tAMkcxrbexKLtWc2/
7odCnB4K5k0bgHNlnBDFqslp5dCNgopwCM5IdLazCaqPNVNfpWqLGrdxIQtFxs80DgeCEQ27eZe6
R/5dZ0GM8ndMPqaW3uo/J88XkFzEErYDciYl36pDq4TLpHNNo80uXpTEbChv72sjr6dMIK0FPDdh
elR5soN2hR7d5y7dc2NlWd6KX2gbec7QeKSugknjRyw2Z0pzvip9Rq8MMCTcBF9CIw9+rFYraYmf
dELHvV8Vu4cO+D0NrwmfEHkuhROl5s6smi7UqU9Z4s2ApX7JUhd8SuoUHKgL0YKwODdfy2aae2K1
JHvfV/waUTlyZYCoiXNxmrmeetb4jPb5mGcIjTPGU4RpRvXyuS5q+V//bEA7vslbSxRafQdGCb8S
yFa/x+3nZO7btcVuruKJoZJ62e2MziSnSMxeRCciG+5skebS+Fe+M1fFkzEpSq0Vqt3LmFZyBsgt
TdoC9vgUa2Bo8m7+dkjfaR96ufwE+k1+wRdu25UKxv4iFIXivviyaSZFsXHCQVp257yZ+o3oGyiO
Qm6dlKyUzTJTUIrFAGxxRO/KDg7OLYFqNfnOmyquMNyCY5gmG+UPiLkB59FKWmXY8vry2bi/jkzl
wgA68UXsxlUBctYGs3q8puRXDPIQXi5TccuLi6TzwYBzuHuuReU6oNRyn1QUjFvXPPssVk4TobMX
Wyzb2WXVu76cYVrEzn0nNwTj8l7+5p1i4FGYroQNe0pETBeVQ6pQS8vdpUpNyAUrgVEHr9xRfsTm
E45sqLqRvkeoByvk6Iqfswn0TkZJOSpC2c3u36GKW8jDoy8Y79LzUeynNdoPZZ0aE8ZPVjEFySXr
96PQoOYb7bnoSkts6JJMU4OOLnaNrykxA+Ni1fmDj+j2VKGi6vSWutZn0qqKhfv6fQOrhnTxhc8+
ctQPrVHKAJ3frXZLbhYUNcJvuLyNBXeP2twVOY3jVuqgASSt4SxzbJZ6PGY0pSp4B7f3HepxEHgd
OXQOwCEMw/4Tuzto/gBSipQN7KaolT5Ejm22RrYIxNwwK8pkYn57+RiV5Jfk+K9Npn2sop0IIOsZ
5u8Yje19l+tURdz6Y/kLklZaoM/PUzmJ98M97Ey6TpbwSx2gbe4iCTnGAd8KhVEWhP5q1mtUArrh
9T4kiPUW9BJ6MGVjGKCfNqNqO5LijyOaD+gF/tvbZKxFq3FJGxLCrXawzf06/7PFd5TSnufctHvG
gkG3AhzlcCX8lyKwkFzp+ga3b+rddDavJhVO9HywbWQFAssTBEYm7mGvJYaGAg51qVXChaVocUlb
f37ZedrvzO/EVWlX2hEI/NExRYLkOlhE+/V5NP2OC0yaQmyiYITcenp7EZsCggm0yWxSQeXuo3OM
lvS92YRp+CocA46HOxkYPNlHT/a9vTb4J10dRQbLH4dhkyzhAMf6Ru76RR2u8Bain2dpIPZVjSZm
4rod8otL2ZsOx5WwPf2KACIRubmPOqapIATlrWDrCSbJH3j8/Si2Q4iXhmAbyERxn0Qbpxgd2Jsm
+YYKwjvzt2YwGVnuvsU6A10Erfwh3XhqL980mWYNmLemXH6FaT58j1pYmhcj52ZnAycDnW6ugvMU
v9zkf3DrpuNKmTTu/u0X6s4rj/NOUU2cEDzxdn6woYtpYzP7YPq99piQk1W6ejwsVDdiJc5D6RJM
x2v7lw7JCHTjmJf+v6WieQxV+lqBuHMf5Hj/VHm1UycInhIqb9ENvvEjx7i69oSotHfSBbpwenkp
IyeNk2MPvtj9dzEuuCWA9rnv8BAlIJRsskz+TVmHkF7Y4ZBFaEAkl1yj+SGnOCu3PcSyp96MFFqN
0cDruQ7wWgHdSxbbIGHrrM0Vu6SS5ILXXjO9tSvefN27nweE7fRMyH2JMfuJqc/C9gRgrXG6heJ6
sTugnldUq1M8DPR1r23bcTo8k9CrcUE4/kTtHUSpEzy83+EFZluxWjHmwJS+qcstdkCOiKiuRwDP
YXqz1U7IsyCitzbgMvuw7/Vq8E+G2kxce9wePicvBdP+ccN0uDMANB8Lf8s7657dSqXlIMFvi09Q
+7qLqwGt5pUOk34JTBQCVYvwKmGKesd7Kv4g5kAC8/JnXy4vK6gTJ3hGjxBh0m086yX+eGHscOLz
V3GMUW96zC29jQuHn3C/0zoT5Ia/LX7b+KHfjQX8Tr2AK66n2KDQxl/vY9yKpjcreI24uISH99ZS
j98D56mdBvlyYEPIF8wS/UeH8/eTXJYunGXjdnBd3BpVdEPsarrsJzx/ic+te+2sDGKIKske0sTg
FAHtUlbZNzkdgXK0Cr73xklSDCXBH9T3y1Yd/fltqESofAzYIRGgiNMbJdjmn2VPvIQz/fIuoYJ/
+CqHPl6qT7AUV14yzRy7M1GZ6WdLJrApXW4q+ZmjQmUYw8LuQ4cTI2Odv04/7MgxLsoSOn5SNKP/
IAexGwJ21iZuGeA92ReTuUaRH5fEh2ax65QFgCuw2OFJC2/Xa0GqXldiS0UKDGMSJOJvlJ4N9+iV
VJYML9Tq/3wi9lueCL9+rIkJAmoI523d0AIOMLYJADK9xpJSvlO4VSalK5wikEl8XLgknUaBYIxN
cU1E5M7ykEZfUn6JXFStre7Wr/tx3E650JdN+koY8xw3+TH5zqJkOLwSaQS6CvhI1CuOM60YtU6Y
2v6PJJzv6JTWEbnUnUjXLHAHE2DwdigmCj4nTxzuQNFZR7ZXRqUoKMC2+Uez1nh1dN88ovkf8M8j
WxlEYhCJQlG0dKzbfnFN2zfGusW3uTMV0dDkAYaXoG2i7ZQzfUDL8urqvxjSlYKFn5vW386LHvAu
6E0T1gadvJxZjkydaxcP/Ro5/9W4kp7q3lEOqTDGThEh+KU5CvWqVjCK5SNUKu4Sm96pL54HE2LN
kIbUFQKjkh9KmjROXwotE3Mhkgf5QrhewFIMU6gPnH/doRl6qTYwmQ+SFuWFQaomHQOdM/5+reqd
ZR99aqSy4jZx5ipDYQI37q5XsIiQFsTYgvKqrl9rgU0IdhUq1AamwM4y9F6Sx9rHSMrznjrCicDb
kVA+ebKbxgU3Nw9V2Z+AuWSw3uzl++GueQ9B/6Fb5ar3LpD5MdRA0kVHfZcAQjShUO6hSba6ThVj
TKLHM7SMf2hr8YzZ8mdK82vyIUept5eLkRNEYHHZdoyFJwQ3ksD6KMl5TLiuD/Iul19PTjVZquGS
uwrjKYqaqJmpAxfAVwG9XK98O6yKW5cIOczbEaONboHH/pUztP5WgVJMIGtYWQc/vsoP5PX0es3x
Aub4zXaXUok4Mq5J4YfGtpExj5pwcH8mGx3Io6oPdxG1zwmNqXQVajzv49ST99Q6Al9qJ266husD
YJzhyI6F9LmTWYrUFke803AJscdazxz70mampWPP9Pkrnrd0NvFxZP7V+oGfGh28+om/+PYvRUOk
/6jqAp+iyzpa6bV/C/ILpYx8PTHvp/IlPEUuj53d4CEQNqki8S8H1lq+HRXHYAwpwGwms2K8UnpZ
c6gseXg3EqhsM4MTrFdJaJO0uFDgtzBck4ETVCErXcdMor0rRvwq7FHPCWdYxif2dT2k4nGaTbkg
7zSJF75W99PZtmgp8Ikimz93he6jV5kmNfG2wMKTDvOQcxk/9Qu/VYE2D9Zczkls4koqNOrMepHd
jADM7E5DW8B/b3ehrQvg9Bco2dqbzVbvr4IQaRZeK77P+HFEh+dJUdfnqQ25gcuI7J9RAqJhP0I6
HZMCh7FzuGpJvR5J7tBoN4An5p2ZeoiI64vnJM0ZLg+G9VinIuqcghrZtJ/qJsiymA8L9vi+CMrP
677WnlsVyzRUqHQW5iqwwSjG2jahJ/u7lPqtQga6ZtknSAKKarbbegF2TBtrpDBCHzquKGS1HUiT
5RgbbHgruONUeOR33RAnIKRrpNgJG+MQPQ46/+ujo0Pw+XAhBlM1bDLULN9zCzFh4Pefq0/jswLA
WuOEwugcWJ6pI7XHnhdo7gfb3G5XVinEN+1ArSIKSKKrXmm2mJ1Ove4oI+wTFRHEUkVvsUiRYiKt
WSuNBYJknEWAmpglvBIh1g37AnaQHrjHLgy9FiRDF1t96O7ObyYkCcmSGFqfArVK1cg+ixjnxSC1
6zQekDH6W+DYZGW5aqop38mkabfLtQ1pPuYrLh7zeicYhvwBFN8M3qUBzS4S2ut4YSjxCSFWbDVe
GLAaTQBypUKo41+JW+/FLheJAym1FuFYIux4k4fAABfVQoMFK6XJolukB2jDk9Hp0vKsoBh6AnDk
bN50yKMwNefCijAptXp+PAs3LRq8NxcVzzkpQttuRdTBaCxXYUbCsE1v48IgG6VWq4e2xhMgakoz
60fdwSoDzPQ6guz4BjeXH8NU6lsfEhpSK+2nyEnJlClDU+O7P/rmCldOjcEDYbqR6/BZ0s+XfCmA
UXKF6Qn3UMD+aH+SPLxWl4q/s9lygWM9Bff8HYYM08ZUFfpmLEYj755ZZ0Ub3+mrazVMqPMFTduS
VetTGc9/IVQpXUeNjUe3emeDxA3rZY5gnWRrbo2vtaoESm4jWjLV9fH8Ie7zxU7B3XkCGHIkhUIl
gyhV30rSltQfJlEC2cKUCClJy4SEqxaZNYpJKIdu+o2M04//AR6Y2AATKzN0yloZOe9IcMhHukaA
Zg5OeptQCry8BIeaImyMoNVHjcx7FHM9Sn1gx98BLbblC0mbKFIBLqsgvEVivb+gz7DCH4XbDbuk
aCui9mQDPJqvc/rSJdgCclb5FVkpdUtFINuYaNjQqpPfnxEQmRCc/+SM2kLnp6iFNaenJyskGFSg
wnJPF3gzCd7XB7aGXU/koaV7Z/kVSKPh75RPCaIsz5Eq3xFGRmQLGt40FRFQIYqzT0AgNSVRG/Va
EVbOrQbJ7do88/jV2ZkEmeo5p9vUZzBzdba4kq5jlvM+O/PnJ0y621TzT6WmjjVIDDfLwHlrpA24
8hb2Jv2WA4Z0jSYAUgl3OpKWvXvNDvyamjAKPeYpdtASR1d1K8Q1m5Nn/zDxRiWonVaVuQQrMW2u
FZ8KEkYyhz5KHzxSpSllHfKcq2+RxwkQmS47oyjFRyfLkQLDnfUVSvEG+CkSQGT0llTpQqJxPBRT
NNNQfRlIJZsemAnz0QruKhJmoDuiosNtSBsWwmMEdQoceyP7wtwXxNIOnXxQuqWWOUfkLiqzA9+C
uB0WIYupL8Sua5oVoAlyn8OPbMeOgUtnB8zNXxb9cQGpJT+8FbGfdAroVzv751wh5Gl0HxpFA5hU
sF9mW673CeL7HFphbd+cwWbVTbrNnegHSSU3/4jXpgg9+rC6AdRwrrwFr10zxuqmN+okDd1iXuON
WKfm8qmGWMbjQlg4mzfyvzztu9FQ/snyxH538/BtJW8QQ6MnFEr3jB5bgTX8gYyRfdKAWr9eOLYE
b8ng0k6puTe3IcQLDPtlrC6MyTp8tXu82oGrNqSGXrjAO4jj2tSkrmsuDv/EP7a6vxP0GD/eWHZe
XMNfwBH/mG7wzuA+xJsUcXtuoTRSCC99U33/t1C3sS9hL1x5M5GDh6cyAZzfq3PvIBSefi2IeItV
yGhTKg7aN7gbOPnY780FkuSeS7KbZYEmhSJscj8Wie67fgC1KEhaLgvD0HlVnYa1odbg+Oj/jlmC
5WTmLCeI2DgxHKBnsKIXt/3hvg/f6XZlicHuPVgnldZNUuxn4Nd9UWQYynxTBvYiNu8jMfeUvSsy
xqC8utE9UDrszwYPrj1RofFkFU2q0M+vXZd6JufjQmii80b+PpoyqCDIvglkF/svtIrof00Vwfcj
bMZE+PvJVtwQAF/8r4GdpBVuyFeWPf3NTQCUWuokPncyxcgh09xJmN4QXzsyHBWnM9IlkwBcaF6w
t2Qf66NAEQGoqXrVUu+fjOvEj+QnL2uruRFkwx8PhVBFRjRZK4oqr7lVxYPkSGm8XtmNA+G2xU0n
8JaNMJ1brvrVgbCI7I7JJlbYIo6klraESz4gzMBu248QwLZZ7ifroxIOyg82ZTN++7TV+5yorQ7V
azyr1YS+MuofjAAyfNWGn/M1DiUQiSxAgiF41Gs8F7duyMk7LTpU4pG9skXHycnALW8UqYAN8RFu
S3F0JBvbVuXSbW8hXAULoWrHOdBizfqjwHrZAXq9M8v8pFlo2ajVtjno9PAmnjuQ3liw2NV1o9cg
ktACODeFic22zt6qmnOoD9PGVSeSJJC3GL0QJUj7tzkupNCY8m7bbEfStj5A/ZbSU5Yb3LrE3He4
v50nnGwjjW3WvsOh9Sn4FdCSVdSNDzBl8Z8uYPsjv6QeVIUl6zqUOFlf7dHlezaS9MzoomPopU2a
fIMF3vmELxdSigndJSySuOns99VF2JacebrSad2R24/2yAghlSTgbsj11fsJO5oy1d2iBC9z6XNG
IaKrSJPtLe2+IulwGeVBbOZg9NznpEtIyF8qIOk+cz+xBnWtnqBVf/xq1jATVUvx4Y/tp7/9sHj7
+u2kfydssRjhV7IwHfIuqO9xIyoMNAh5YUjAPS3tSeWqDVQ5TrZbfZVclw8kNIsq+Lpiixty6pD9
d/xKmcYmJOHQJ13hAneM73gnbrvX18bP3n/xCuLCUMLI3RM1QtC821Qsy+pkJtFr8kxAFqs7kcxS
ztqac+5clOVn1iMVGLzEm6yRTXcSlvcV+ucmhNgH5UhmuOBU/U6CPki9lMskpefLQYOoY/y8NhPt
he99UmTmtiePRPsraZxRzS9o5Rxv9embGAPTtfV2cEfINiCmhDBUntdx38KQoR0H4nMzztwAI+l5
vl2VaEo89cltl8kdKSgc4CiClUR+V657us1elK/3ij1xBwRpMjEct0R+mPdkVtZseAGlxUNKUyYO
9/Jq8xZ4f7pESUVjqc6GjwKnC5HbNdCkNFkaIgHbButt8a8t7Gr0TqolDDLdcL6LcRw/PMkrazKa
IPeM8Dh+DjoVlUuewvO/ofsord9qTYrZc2LbVmPsKG7ZWo3FnHWAPgB3H+ByHjDZHXAw7Wg5z70l
th8bnXCydW21xrYQz7cfknsfoRYXPAR1oY4gXffxWjfo5X2/kvZX4MNQIj5CX7HE11sj3pCVsaAl
CXMD3wvFtJA+YtkWgdQfH9sq8RxJ913ff6j6LA5fmRmt23TimIleF0I+OOwCiUmyx8eudIfyKjxW
b/MgWg0VC8kz97tUTWaP0pjESaLFNqJKMPgFSeCaaILXabbLfKtUFRxi8W2zDKJ/ABKn0VOxY/ki
m6G3a7B4It7q84zyQhIdW37gXh0RAerywS9xJAmdR/TDBgoRpbFrwtWMnQRvcIskcwy9vpBgZ2Jj
Kn9THXLvFr4O5S4To4B+dim4DUWhnanTjJ8fbHVRLnJIbeTgROSw/Di6mP/oCEAHadWafLRmy5SH
y1UG+he+Lbx3gavhoubUNCQw0bV9L89Jsnz5y/KjoabpJTCU9r1Fgmd8pXTDUroe/eKMmRxUM/MJ
6MPgfE1cw0ki81nqTyiYJtAe16Go18W/TMuY9FGvnSwky1ar9H11MZeFRNFLlX4Yj902NRNGheIR
Hb6yiFFJT4lH7o+TKgNW9nyMXiCtyohQNmTWRNlgxU6JMb1z74JoYF+eTITKH2Uc91PsdVor5INn
hUIxxZnLtRnc8QacNM/BvXrgMyGoE+32zQIAI38BWHrvoYXUi9a4jCt5iDtJIFC51wNO+9/wlC/S
Nwzfscrh7ZAs3J4ApKcrd1/2RdIvcPk7E9t9c/w090kHUw4SsRbBhjOaCsj4RWJc3d8yVJSi/9Zj
zSoX2pLOCZA9nQp0ITJFI4fGaQAaHK4NGM6UHuOWjBsSrV9+rFHXo2jcj2aqvWn62pXQwMxvpbo+
JeWFiB+YZ9fDy6gG8ZqWfRaaCOW5lYHxacLM9LbljB7Oz5JHXzKI33DhcAveNrd62LAfgIA0i0/a
AVQZyIPpPeOy5sXDJgQvQA8PUDAJwepsv9g+8UqO6K5dhOti8V61WRS6fb/vxn8PjkazBeI6LpRw
ikiRyTkF3Xs+d8kolI6+uzpl9bKeBLiLJtPQEvGryr8CKF5N6pFLIi9GK7xS/1iJOrJNOL4Lw9at
PMqht2mL5wcdEXVNMPR4v09m4ypmRAZc9RW3OARY+y0MRvsPSabVouX569eWYHJ88vkEg8/hM7Xs
8ptf7jSP2sDSHS2eV941p9/u6VAAJBT2By32Xis32vVWgziOvX2AbaLB/jWqe1iaZ+vfp3Y9ZhHT
wFGCUagQX+PFirrNeFk3PUDn4BnD0floJ9W8alj7AMZwKCEol6+lqD017ys8Vesggq6HB1wIAJrq
rX7L4XPFPIRmQpUuhBv0Vev5dB4EQUcYe8SIGrbe09pI49PjnC8OmeXEs0q1S5JR7Nq1R7mbfIQd
+p4gS3YWppFGenWLs9BYmuxT9zcIJMQsKT/shjRZNiwFSlfHVpAPj/TtQ2r5/iCMj+TBW2io++Sg
hBHpZqdc0851KUScfTc56C5dtzYbcOB8T9jTgsQQkqlwCUbCLnYpRlShawMomx8CqPnETEUn5A4U
vOHe3Dt2706FsKJ/037heohixXR5Iq73MLL+osALc7LXUxVsZxMxyKghT6WOpM0pSdlkdzUnKkNl
nbQyYX4EWj7HuVZK0z9Sz5rHDd6cyX+sq4DRnOaB/nT/wcj0keLFQbI9L0DSDAmwQWSa87lJyhsx
TvT2taNwVy9fM3raLqj3xaOx27wn40oebH1ENmzwy2KwdeF/hkuBfy71kg3NvgjoXwzsioyE2o5c
sFxjcWeF9RZ562zIhjAZAF3KBtOYZTmIPiRmDF/1dUY627Jjg3+jCO+OEiJ+gqZS7n6nNybzy+6h
DOjCVsnIuPhKOD2WB/5YUf6KSZu8K3xw1r2ODldaDEFFmxIkRGCjBYWbt1ZAT8ecDhNIZ8SSsH3Q
ysvW/2mqptQukU2AuJvbREIg3LbpNlU25GFmUYF/p3dm5rBAs3qeoZS3cemtzumYHnINHi7MGMHk
lX6bXl4NX4KuufB5Rjt2aFCzPUAmlxlp+cVZwlwdGBfhV9fwyQ76+zqiYKKpVufTDS+raKcjV9wN
sIqeTLGc/G6j7O45hWYVuJwU310+34Pd+sOnfHBBlDHzyuFJ0/r4R4Ua72j0hQqAacGu9gQzheWC
r6Z3DkjSGOF97ZcbP0R3lEc1+nmOD6noQG3ZF7ubXnSokYG6RNM6XM89JWks5JC99366gzOypsIX
IPQG0w2NvbofiVjhtbNNciFEVbyc9C8GJSe/PVtwqPtMXDiEdTH0zHeJovKYBIArkjYm0c1GFooA
wEQ4tvoBFT4GiCc/iwJA2oBQJHHsMxxIb7UKvLHmv+bCBjeH+sc5SZjJBQCDngpdTtVT9+LpxT9P
UHzk+OaVkzaSW/mesRHOqjwGPkk1py+FGfBFpiVClFoHXQXQMTjIGWUzI89BXKXsTXxE2vBxAwss
BWtqFZwQb8kaOGy3++2npRbBsZGlMsTM/GcO3w1RO3xBUaPBaV2TISufXPVNVcE2HkUGeFprrPdP
3vBg41AYP536SWu4GBbpwtJbZjhFVXbLD0kK3bL76flukIBPcsQd0yfo7P7r1J13Gjru0x5EKUS4
z3aQoobz/RiNBGWRhAc+j4bwZQSjKMl28X7SzwRryKhAwbPINc1ljg6u/kzZNoIKOIlGqKyKH+JO
DVXVS5C1xrqkrjS1Az2gHN4+tsL3q9aOtNBhD2jjKOntRBEaVW8/Z7VpP/Q6Z+uaOKMqxoKKXiYZ
PK13FUgDGqINVs0xwoUMyW+nYB2zwHJBokWek68QXYUb+hoRxnt1Q+F0ZS3pt4MxQNW1LhZqumFw
bLXFw33w8tFuT38bSim5xH9hQWdUJRzL32hcoHC2WOlGMJFlp+F2SD3T/UUdxv7+CCs3B1RXoJZb
+qa9DE2q6nBc6TmVKhKIAGj7iF4e5ppHxAOSOxFytl9q3Zc9WuvhDxGv8ibCP9zM/orMlRBCXUiF
QQ662cE1qUf28lRqChUd4WZI3WRNz+VvXUYatAMbKAznTauwuqpjcRbIR8rCXOF9Qn+QTnEjC6EF
4mt0MuZtR9Ec3IBTi6Jpb3hlUgBtTcjU8ZZCttGA7/Nhrz0yEDunRySlVmOwpF6pQj51zzjLBoEw
Nc5I2h8FJ2HCBq1mXj6Znjx1yiRBgZePTbr8ElrrvHrBHbfhGTo6TQW621+QhZblH4hj7TMGi/om
MrznJRR3OcBJv5c90GlwmFxQZIOgOzYQt0M49Hxr3XX/zyi8mOO+8J17nTvxohY2Sdt4h5JeL+9R
brr5Hh1Xr/G/ZLGKfVoOSw2nNyijVlvfAhNYksN9kuOtWraUusBVUnu/PpN/ueT0YAHghbmNHSSS
rF2pvF9o4wzHkzWwZF//FE0dB9DV+zhakpKx5GvSyw4v6DJTJ+jz82l9mfhdFHr4rEI5FanGzZxq
vcKCWWGtwBgKYSaRvulbH8uL0kvgaJhaszLqepN+jp3/qPHlc76ymARZSd4V95ezNi6s0nxFWEbo
ktLCkJKO7U7OGj7FhG++onKAwPD7EKmbxWu4pmHIiBcBuer9U06UzrIm079z6FYp6IYH/oeYAzny
3vGOwh72E2XNavoObE1qZUg4MbzkCyklhUuXMHH9ygg8/iTWp79qr3+uxCQgKj7extfJUQkX7i8g
SyUIPuDf8IS+v8Og6RuTSIY/d6kJA8v5VVS5Dh0POGqa6VcFdq4uP8sGbA5sE6NAdtqWpq1SJ0XF
TgeWfSwLfJKrKbesd0DsgE5hqDY/vFjLnINKuJI0xH0YCo5B2/ar4QeZOJHK0chjK4JCp7b9XO5L
shFGRGOONhxALzpxoXAM4w0hy5gxjEuFeytfsiE396U2aAcnvWzptaWpyJB3VP4hef9oQeLOQuKe
oFlpi2sPiMVZZk4nnlDzGeu00zHOgm6JnDIwb/HcMwe0ob6HWCgk1zYdv+o4pwcM7woDTjiiaN6j
+nW99YBYfwV9g8nN/047DB9I1yuwsh9zNWOuOSJsBXX8ujqhU20ZSLpv2Oi++nFSZ+nANCwuGvwS
cgg8l08+pKqowhj4kShlJ3T4JWL6UtjIyCk5HkbqZzwm/S9mO5YEC4bYXw3Gpcr6doqkPSE98s/H
1MUo2qTNW6oJMFudqV5AudiOHlKTxA22PqywmpsIfND7sOxPSsw6W4lotfmMwko0oCtfEdVHvcPf
d22Rx5wZp1+ffkpfe0IxkGm7jp3dleNG1qkJAJYWgHi7FlyvvTsZfHcehRMpv103Z6riB2DN5WN7
h+6L4Bifjcom3nV8n5ZeMGOZrHh8z9QskHHjFQpKkznjCQ7hxcKGCARRGRNr4dMbpge7Mo9dCV6s
t9dCoFjTpUfj5/cAHYhmIpqn2UDG9Smn5tQ1+bzftkxvHQLJr+YS3YE+w651/3En+6q7bAHGe05U
6OUH/HL4TA3Khaa9pCalEr+srwgiPrkjqWDi1OwI6OA2lb6GSpOGvAgc1e6RA9dd0NA91VbSr0l8
/iS3OtOjvPzLInDX/jdJogIcww3jmmMUlcv2oppOqwvYgW+SfhyTIcszJVgdPmU3VoltyQc6C4C0
DTDv8StoH/0oIKjkkIcSD6A8gdVSnF+IwM00y40aIZx3/IQs/vfYR3rmyPT6ssLwBtZS7uut+YS+
FQslpNuUnrTXh8DpdlBoCuChO8B4MHb8W7KvGow/IHW+lNuuR8CNQT2N9nEMfTUecsf3xOs8X8xx
PlBeK86uRMPQRenTzsuNWOqQUxoMkZQ+cdx8OYfJmQ/Pt+dD4xMUiRitmWrvn7bht7qkZ13yX7x5
kBFbrBZSob5ChipopY2/ILlYNT6lMUawUc1qnwhbmDNTlnz3A+Vmt7Hl7Xs+L2ybEW7EH+ccZC6s
qvHNgmkeKmBKVdUl52PV/VLGE7S/Bd0iAj9rKLwZmFQsyMTwx618Nep6dJgcjSW+B7WubXM9HH+R
GBUZ91R5rEGFhZiHBnAu4pLQL6Wced6+gI4TAm3ZIymnZreioX19mJ6CMEhR3nbNOYa+gRlvtvnE
1RvaIP9yCUGUtnOgz3z/HUtYhIr688iuTZ15bprnzHiQgZIaPj6On7p6RWBSDXO5PPHdISvgUNzU
WCgVxiXhHxeLNT+C8NphVQsycIEQFKYgi5o5HAnJHbsPka+p1OvKlT1ygOP8cBiBTPbDcEf8Gi7u
8XfS5nNMM9Ab5m6Hh1uu15dEYOEQJC+7Kpn6yXRnV+1JjDp/B2V2LRIMY4EnXVdT/0aJ+99PwH2I
g3YuDJBuDjFZC0joFNdtAhQMFH8veqko1lMeDNGa+0uOJ0Tx9F/+tFO0pah/nYDf580cOXVLZHjF
9efrM+3g2eMsWB/8a4GzRYwHzo01lBFjPlQAl/YSFCJU6Ce+rOoWzCBO5WVxeNl+sUKWA55mSm0X
Zq12AZe2whIwSFIyKubiGqI6dh0cayonVS39LYVZ/VH6NZh4fHKWP+sIJ8zla0FfhCUfs6e73zut
p7dsHG7vqC9/l3arSKlYLqdgeYE3g9ZDzNu4pFZe7ZeMDegbpdyA28X1AYmB/FL1k1HImxfH34Gh
8CT0a9Utnc8TNpkxNMiD8y8mfzCL8t35rQL+uUBXlstFWqWn/xq47C0TJY5TCeOTR26rwkpLZZXQ
j4XcEqC/FTGJjUx7Li+TD1NLPUQzKPH8ZTbclZ9SWNhTHYKBUgLZpv3SY10m33taun2WVajAHCLm
pvBbPtsy9dU+i5WCloxhmZPKV3aW1H6yktngbmCdjUfRawzIw4u/HkqE2iZ+mE5x92DdnNrkfSER
1y4z+d1yRinuvVjvmxQJq4sf5o3pVmFHjHK4C8XpB7dQ0j6q9pW3CIRK5D2m6W8NfOEGyETRZZke
CNEFWKI/YnYLeVa5dW+zpLZg4dZddKcvMv2NGcw5D1lVFwMumy6KMbfbdT+JzktHiTudPSGQphDW
/AGbWccXY+f6ZnjNiMxEsRPAxpgyHy/LfNnpTZyeQ6jSdKCzgO8H9RgmjhuxMyfQnFDSgysXj2zg
YPtuviPThTtlOSqUaTDMdjFU6yztlDnA9xQtNuUQAyLP1kWQabojrjF+kMA46OVOZJdz722SO8aY
yZYkj25f1l15tAgIh/1aIg4C44DmX4rYJthdRDHSwjr4nturyqF76A2Yrjqal1Dbk8vnSKZoMpNn
rqRePyhgv+rrJC0M8kK61D54iL3+YiK9XH51bsnVek6N3yh1HnoacLVXzrYe63f7Zrzt6qB5ZkPY
75I+HGbpipdL3R+5iN0tRWbmKpbJwZ3zt1QV1sHUETzTGdCBIenAcz+yaCDbz4pHN39H3Li074Es
GY2uI+I1h1oOUcIBTzEu5hw0YVRXzPAh8aPJmxz4+kgxL3iVcCZjFeTg0wWHNEyn/oOlxoiUFytv
iBUu5ig2Cm9Ge0jHVpxPXSlSuNV+ou9F2skZ8tlk5bQYXL40GH9I8oqP0IGE0v3czkgbBrebCuqa
o1wQrnPfBJpzumrqCdEe0CC8MMnwRkDJd7xlryS4+zTaXhqTCtWxMCeAdoU/g6KE21jpeI2qikqG
TnQtflgJ9B0NtJkCdE37S4OGgyHRxUN+hYDsilqRpH1sIlCeLINm7jg+tCrn+cFnNN/UlL/HiVpC
W4B8HP+S2CwEIeCP/4t2vlvP74csG08n+iZwpKf6QpuzpoR1FlKbWcOKj4+t9NPGxxnI1fEfQzL1
pHnwqdUaHy3hd2n5ACQ0cda12XfDLUCWCXbfyFy8uqTbv7RWwE7BEjP2G+sqHg4VbKlvQysWzieG
DjA7Jo+i3GdgdBsu0cl6hF3gLIDIn4bjodE01PWRyTLJ5i4A6pLUrfjM2ii7wjdIWnzQ3uTPn1mE
UX7vnQ8Kv+q1G8Xy30ILsyV75IYbKE5DHIQrCD7eomN7UWBQBzIIx64iOl+bY7mYd8L4LYPdyZPE
3Hgs7e49TjhxOWQVrgOL2RNAZiIfbs8jrVT+qqzA1BvhcYtKrIAekmzB8IqtVAHzkX/7ty8Gp79d
glEiAeMhV/is6UbXUtBH64qwtkVZAABNj3z2gm5+y7ObKrODhH4AKHzbTjFaMUbuGk4noNJvYsLk
B6WW8fLzJ1a/yYUVzS6yuS+Oi8Gqiwj91GjXPQoN4tSAvDUiPIfGD/vUoym3IMk4ZWbBK9BKkRmG
Evabz84iNANBbmXVcs8TDwCtvJzkz+yUMwClsWGVYABmZG7Zvqpt9M6w4e2lYecogNv5hsb5GBZS
MvK5eSzIITi+9lDZ1WsAOrN/SjNGgor/ZHVbE00cVooIFZeuuDZRI1/kCDRyIAU1XeRmr0o2tmX8
Sj0ezhCPwvzJi1NPyO1XFjVj0PdB9QjUvS91AWGtPnbeash0UM9tNjT/NvhWLr8GunM3wWvhj4qO
VM864bihrfYvDEEt1MWu480LHumZcD55Zq0KsREZUWMVi9JMUjH9mNcxmBMTXevmXDA56+3kbZfI
8NjWFkbNggmUKwB6qzhjIq8oPWK5uoqehEFeAGyL/LLF5eAWzBRSWCWL3D4vaCPr8YLkNz+B26wj
ywypb2/RTKnvGaO23PkrkT28SoZbWOm5WfzBaf8NWpgYhkjjO/o6lnQAYcKhVTjHQ7trKGLhJ//Q
hA8IEp6p6bg6K2+Os6lROrX25MDz6D3b6X381+nhKmK69Ky4OCVnyKtAg1jLtI0p3ZYy+DPVBXKZ
9RN8m791deIQM4GbXq6yIxgLIZ84gHuEEyuu8csRHUhBEfe3nxp3ArYgskLDPb6J/QbhafCmXBfs
QOs8OkyZgmoyLGyJkFk+2DVgLqq1tTILBC0vrD1BrDyob0UbCKydcg8sINN62BcIGmXOsaMQ9zln
Tth6iQf1JsmJltQUW9xsOAHPTsAKFOfz8zxYXYLTM0GsRm6ql3MJwzkWNHE8KroKiIcoVmOiUDo6
IXrDXjQVXTHtfu6aCJCjbQAZw+Y1tMI9Dc7Rq6gBhgL9u48pqx02PMjvIW4E3wsAO/QTdTu6ELlU
McienSyUpFVX1hkSHcqzHDLKqqKfVqpDl4FeRTZRm3vXzsh1KyStsdVxeenkF6GUZgGQJU/wulMH
nOrJb3gdD2hEg1ElE7c4gfYEBn9ZJzUdz0u+5we9edmlxE9oLnw/QXG28L9iOY2SmDx2qlW3Fz/6
qiVEIp7CPRp+EplGZzQHWB/1rMOll7A1cQezZ/uclKxcCI3QnHcI4i0msoR177AD0Q04OL19U8Sq
ZIQXHou1XHc7PvtDSP78HVEyIlBBv5rcW/7Dy4IEZDh+UMyJ08EDYPa2X6uBYJ54cGeqpNKb2h/I
18R2UQaQoBcXgJlttYwWY5IVJnTm0TbcakPyOc+EjaBqezkPY98Asv1va/nMDZfgOi7fvR7RQDMf
ccYibYWvx+hlBpW+iRVSS79vKT1J5MCX+GRlqJTbmNTsvmb5R5tGCG4Zh5POWbECHsBmEgYGvqhk
+YdVgsIBisvwfMtf4hepsYVUTkp0kZ/AA/uvlz/DKMErDYwLNnJAdaO9V2Gwsz8QuzYGKopKA7WY
N1Tp/VFBVeCZ1pJyfy3ePm133K8DCAxnMgydk5PINlna4lEWTe/JDICTUSrSUONF5st5+MMTX+4m
y8BR5GjpDJJQ2GLyOR/xPlzlCOQK/f8DGtWAjpjPFY3pjYL6anq4LwlJCCq+2QbwQn/xwg/AQfG1
H85I4g1s0h2sjBKdaASlRHNHY4W3jOhCNj1WjpaPkVdPqxlGkomoB5iWpY/b2aurbL3Gl2SxGXdg
wNcDwv+YzULvL2IhfHc3+vUIwuIXfK588HzdwnODCFaK/RBkOks9KCFc4H2+LPD96Qj4+ZaOnRbb
0lCn7X9H+xi48W4bubd2OGqPkC76xprRWW/Ys0rf/u3Eqdyb4RqBucuXWm8yWYzMsKfe+zixUjGa
su8TP4CPjoSWiE3SInv5xGizvorEU1T0lu09+u5bIzCGFiV9YlTOANrKNArTVBXCRJRQqjVjwHFw
zEbrk8EnTTCB5E+/JHSSHXbZQUvKBqZsahDcynigMMZm6nD5xpr7AnTSGc3OVcXUcdQM/EthAfiX
gT0LmsoJBR/cJfH+pYTLC1oHCluoEs5+74YGNqDtxs+wHBN53CuFoWNkbUPdNiVabvExyiWkJB5O
SmtdYmUKBSs4vInshQckuxxjPGJY74zfT/h7J2v9+BcUOrwFOsU60NnqIyUjFjGuNmD1eOBM25hx
hY27XdP8TUqXx8BfIASlLHqYEFf1mvCWKisbnfIQQmcrbkmNGNaaKDGbkKBAAHSV30kmf6G7MBMP
xCTIII0sP5eBLEwPkyeVaTDaWItF8DxF7Uwlhdu2U096qSCMUcAEqvk5kOTuwhGGdT0KgOYbRl8A
l9ZHtqWQXXGMDfGeV1290NN14CZin/zBcRgdzyqiMsPVfLLBbcIAczqgWw93hA6Jdwjv9wWFq3zr
jr6xRESg5WBcPMKVE9fXbteOkbjlHVWcW0c8Mb2sCYnQmwGnmaq2vU9QMZwyZCFYrqbD7xmzxs7+
yfKsvOvZZUozQfUY9xe+OJgC4uMjrm7uZLcZO9K+YWlw8s2DIFNzSgHg+mw31YGlMC2Npa/hOqtt
M6wpSVximp49fJ/6WcvQEYmgApUeU3ONjx728rBmzjKMvu1WMbpaYiy7ayDddV3jt7O2vAXdW6S3
TNdLc0J23MBL2u4ZtEEizPVKl6er0qgyn0EksBsxTcGRSMM3yIVp7ursT439E5aaTMTOCEc4c5bT
5AQ+S2WDrXFdXNEm5fB8Vmk6q0VEA3rbsHkFdQytWGFNb4S1Hm/KXUdpwi6UK+r8dOS1bw3MEm39
7kQXOsvwLmb6dyC8WBrv2k60ondPy+YLO9v7miHRwy7K3JWdHRJTMrn3SGWpYDT5ZMufKEyz+dh/
ct4lTmDn2jjfYtMytsUYoWj27cqDEgp1SI716zz6FH5f4XWY6UxS7i9Mqp6qZmP5lPrTUxzaQ1JR
o8ASqunb9KFBqkwd1AykvTORdf59QLIezVKFVte7vm8oe9KdeZq1iV8sC6/thDRsZmbmOoKBQbtW
bYgiyK5uc+GT7GZe5fGiTQR7+K6GNmDr5zok8cSZ4sEMkpkUN/axrLsguNObT5tbieKQwGEDDvbu
ip9RasNFaYlvRrV8EXrbrALwSeQec1us5vaZgDN5WYqt25VDOLmpVgWnyA42nGpM7/1IlVhHDh1l
LrnDYeDIv6NDDNDYnnZDs0OaoKGyzW5cB5awSQNCPfB58it/M/qCBldCmjoBaJ12N5pQo96/Ilrx
+xbKIXxw23h7SoXycfOwNGueyXXu1tG/gNatodtC6QbnoRRuYto7QnMVqaVtTRQ5LIt/xh1sFIKF
PnuVqsSWUqNdUD4RDMaBXga4u2ZisTTmDG1fZZuN6mb/wuLLqg/Ecx9/gHSHIeC+ZSkB9D/dqsFG
QSa0yDkfO3o5x5yk0gyDiSZLBhRZSARz7XI+tOlCic10r4avb/Dq3lZ7C36NHtbybnWyt3Qvki3w
HWoCITmDZ2rbAGtFDNOXT5dzul54Zitkar3MX6XHCNw3k2dPVueHfZ6VXH8KJKBtxey6M3KuQV9g
Pj9Hk1Y8Nl64zZrUfMe8vM7KyElhACu6OvBZ9pUatLQQkGCqOdTMQIxwVsXf9ZMapG1qtBNQdaIi
jJJEkePVo0r/LJMwDr8J7a31AODwXwyMWFjcofDmIuD49w1LKXe7Norz+o847W4JHFgPew1acD04
O0wB68W5qAVyCsJNCRcKD+tUyA+9eD7mLMPXyPO0YzjyzDV1xI6szX4rG0JTtYe0YMCfWu/up3T+
w987M0jwPvd+c6/M6tX7QfcpRqQzAJTzPu/kCLZmdLho2DnHudrLf69R1S6tNMP4W+U5IuCmVzsb
gtylxaAtSqBqKNeQ0oB08YT/aLsWrwPOjv7JQmTmq9JMW0OVwXuol9gudnVxUySmdVggaf8qwLcV
qCR+xZKwsmNLVYFblHZzM6kkvdjZTt+vWfTfOTCkjpTFdaZInLujPT3vzegKkNqlHGYvP8QrSf5U
KQqzUhCRPSHI9aah6/K5G88/ucxgFq6M9aWxwqC1HjO66XrfiKfmA84pKvztpTw1spcVXcwKkUNK
tdwxgr/yYdiiHPn7G+3QN4e2T0L3Kv3LgEFe4OtzPLmNeepMPHC0DfZEVKXmE2vsn342kc7SD3TS
EWUrGqJw+RFVjuQoVnttS92NW96qBIL+DJLtfpiX/u97tBulN5xzj3lq40cF5T/TJD74LIbuYmuw
F2EXLB1FSDjpSgCrY5Ys+CqVSgqMOCFq63rZE5rzZGvCBFVZtthmbr+q22kHkt/ELi5cVfhwz1+d
Y/ltA3aVXb69DmwZYbMXzcJLa1aVEogjHpChQ23yPIVCzbw2STzLdwOUmlKXzVwueb2N9OkPWmef
klz+oYk+LkZta9rR6fud+TYXhlg1gpMHvoJ+0PWUxhHxbNcXIPiurPs7rkcO94/EKxlSZtJsfn0l
+kP3NIFfXi7PIu2pcrsYOJP1KnJ4N+r3xPmMEVeompxtOKvjBVaj1bSv1J1mSAA/Dk6gt5SYU3tf
bNOSj/m0uW4Dz2qZDzZQAvv54F2NTmjIXG+OH+1l4ukftidVTqgc1tlq+oibIBR88uSzRk0XzCh4
MQDJASWhh0FIeudoqKOp4nwrXcJD35pimmcX65seoRkTqcmZ1yv+O5wxHpc4Oh6rYZXBASQAuBT6
qU5NUG7dTuboqgHZCbeO2P9BA9BHAOwOj+U0NG20JrPN9GEzoIXz7YgHX/Y/GEKlarhQwLA3UQ0a
Gf+I0H3aCcxG+ZTJVjhPpBDDms05qFDJeKeAeqBz9cSMDj+NwPsXumWecD18A2u8kR/P/aqVC0pc
EC4u1yUO39m4+Bd17kkr2mxCvK+WslR7IEfZGcd5a6cMEhuK1/J2apyKeIgc0fP9U6sfbJP671G7
cfPfM34XKJywDDWM6lUSgsgVbvYgQxK+3vRV5HZKZh6aszxATxegk9zdaB/LXh9M+mGz+ffgjh5k
O65drq8G/0xRAWKz8+lNPFhA+Z6tSgtW1JeG3tZw/1GDX8a5CbVt5DSOTh0kWtKRhUmGC6dsk/Fb
QiTY0JwVrAzVwWrxb3JL2ElMMuh/x8uWBJQrQuE85f8Ln2ZlGhpwiwGjg7C6PH6d/uOxGhSSoMjT
EUi+C5fUcUxblMK7DFpbB2IJhXKk1H1V70f+BjLDuHpsr4XfqCe2tbQ7RG+he/nsqQzsjX+PYcLx
fMTRf7+fvKkV1O4gOHLmxa2lCG1CUiP1jz8SQFMEP7vYyU8fD8PMcjbUSSD8vtrg2qT+aKaUbHqB
X59Wq8a+1IO4R1k8IYdCAy0Jn5SVQKWLcL8gnFld9n4ADAfp1CkmCupdzBvXdRUeEbcHGjq5xq5z
DK8ZSreZBv3rr7mMCofRhLRfn5PQiTODxBdYPQK+Uw7iH7L5aVk64VVAkfe81IDNvCtUTGqtOl2d
vjXiD56KTmjLnKvWD75ukFuXc1JzTP3T1vTK0UwDaeSY+KPnFYlnUl0HJ35Lf/lhvqNVEtu1uUXV
WczBFMwp5YqZuwpSZIL6zGeJzCWiFkTVmOvySeNhnpXRohS5GfmPbuUQajlhJIy8yqcd9uAuFdfq
6tIzgfNAIdKfZ5KY37vJVnO4lbgy2mtH/GlVLWKgL+m0gU0QThxVRZDCe083D6Tjat3mG2mhxxtn
OzimzcpNioMypLVuqB6SB0UFBzV56ey9gKQ6Irt60iF6tXTJKAiG/SVQnLod3oM0XfbmstxsWLzd
bOTOUVgbxuqYdwz1nciD/mGXDXRkHaWgLez2Ny5v+HsFag88GPEmNdrhlpGktluJg5d169KF4Zsm
ctwPVIh++YpPkj6uwkCRNjBDLNpKIi7q0d/ZHq18dj5jbKyHeO+FqQOObQ1yqJaYn+bhK/dY/Tdj
BORD66DL2cyLRZXhH6ZF5UoIzJtVhi+tpsDTJKG2hMnUhRSNE+oteQhHzYWZN6ea2VYHQDrg1C+A
YbDHNEI76qRnEF1vfZiNMZlzCJKk1wNQTeFK0qy34YuCocIl35YN96w7kzfPE1x9M9RZBvhHdfNb
BKYicdPMvtnIts1M/itXVrSfwuT3C/umOfccD8sAS7yxwev14j3v9YYqVXXpA5dPNfONND0S2HLN
nnzmX4hxeXSb9VE55GeO1vly4rIr2xKt3IxvB5MtpZEJCIG16Y+xKIr4R6U/OID5YjDCOPjC0Z/e
soGwmDN1rY1he1J/bENnCd/poTQur6WNr84E5dDJN3PfImED/Ih1K8mjj1JWKwVBkoHDbNP3Oeyi
PclIGZoT2oLKcb5dZDtd8ndDJbciJi3kJMKztYX+sPLrSU0glFzpP6yy+4CbUr8N3bcopYD2lfHY
JfwYLuwqAd5rTkb3S89qLCdX39kpkcjag65+0KrzCoaPn4S3ms8h1X5gh5DBlmg69LX5nWzmTQyL
rrswgSkg924YFp4GzV+M0/AJvGYegksOnrVKtdb+FCH2ecOdvBv50NcMfs5967E46NtT8CHWVzOs
tYuY8bXNRPB9pHUTMMcQldNBE5GO2kE2hRM5CdXciIbX1f+VnsmJvYaH2XaiyoWMO2G5Dn1u2WhT
RitEn77y3gFoPO3C/JM7lhBN/v7lN8dP+GjBj2b6vw/11lvshu5oUVcopheZ2uIN7NIo3r1fC4XN
pUxotHnNXbPoJLycndfrnX9fRP+Y8gfp6tEzHtM7qLtNtXvL1I1C1ihRqMYfFFti8PtsqvBneKMx
FijWg6Rw6axLI7fs/DbaCSyuKWIw4e9MacL+OcQ6aCAyllZW9Vyi/TqKBiOBc9CQvOZsOKJgIKN3
BOhX1rdmkucqkluw9BOTD0LYe9vt5P1Hqerq+tyOah+Yai9QlFxIMnH89UMQNkBH/mhSgnuUwfeZ
yDtM6F58Wg5fT15ThiqN/PwKYmwEJGmuYkicPwmNcYvsiPqerfLYoitExim+apqABPEOsCIzyYMH
CpnLhxg4jLqO8dcgalfNGDj0RFB1g2CMQWRgJZex+CPFVqsPF8iuVXow22XSWtb6+FhUlGOd5YZy
iME/EOyVRMYILEfzxhaatVClilT7WQXyfLSTA7at64gqJ5tsN55fnqb9pKCFdm9uN84tzo6T58vh
zttn6UDdGEJoQKebwWhWxi8jN/AGRlY5OxT0kytORFWGkCXhGrJnvkApUME0vcnWY7CFOCbHa4VL
xeZLhll032zcQYInWIf2Av4Fk3yTLtgR2WQ11ZC3b6OFm6WPg6VSxDuuNGa2l3lemn7pu89TEITQ
/QKSnJTe8U8DJgyDrXYIxpkF7a9eILJbCoTuluE+SI6UdSxlDKWjVfb5Jta8+JQ2wtux8suUFuyg
0bekTMqZmaK6RlMPv9HBT7cVS+/nBy9hK/7TBACAQfrsYI1HuVbWhxnpxSlwnzKoR36qbEHWGZuK
/GAXsPFXFOgbxxUIPpWf4+Eipm5Cl9Upi9okbZ29XSimHlpKNUJrub5SyAZl7SW0z396tMoPXWRU
u6P/eCCVjU9eSHCfPDAmJtVuJHUGyVEjt7ZpBcoms0hsXUM8ND0Mn6QOisO1hfsRnB6GKQez+Y3Y
WNoForqNfLnvRnKXj0x4WWG7Kbg4vDYHMpH+uXlnIuBvc07iNWm41jFxBmdepYmWe0i+Gn+IKAka
U1yfFOQDIWOjONilrtu1zz5icL9Mw2LxRGoynAAke2EALERY4Xyzi7so2NW1XCkt4NaIcMx1Eb4l
5DfKeFCZgY0a3gDRWqGelgoH8vWFtoOfyTvBtUIpc+iFYdcrG4b+NG8zhd0SNM3zY6rkEfDrzj+i
5o9Jz9UEGprOUpPuRmmLbFwbsdSj/lWyzsvB+ddVm/ixsneI5ttjWm0j0kjqRirc8NTAVXAaXTML
mU5PwYafXFAN3I3rgxPyliG6H1jzeNy0G9xMn3LE5XrZhzTDEluPYoj+isBsjQ6tbmkPEblxh14U
OW0fD15NuNMdixEMiJYIYKLsttIOtUuZvEpVV2YWGBQER41bNEIu1HNK2CWrhh3Fl7kWhar+Q8VI
fdJbFgtRncMn6IOeA+jzYiJjyzlhFi7C/vpunyu6ZXUEBfwWxmRbMpwJADlM1DFIHdCPEnYGs4Tn
9nwxvYcyn3n+FcrqZfuFyextJ+Bhlbm5ET2omgcprJVhLtouLchQk/jJN+6iE977r/rqBKq1UoGr
wTb5Xrs6DeSskNTzyLGkjVs7MmIg4coPsBrg0GdF2qJSsFk8yiw++ZrMPLNsKpXRL0aMOFQfTwvI
Ww4HszZb7ZORPhpiArurmYkRdJfbBOmAp3KkdlpU/+FIg3BghFgIstibjdOEg+UPofwIz5b70S6d
ZVEHTcBT+1eIeTU8lP87T7KNeRMYMKsIqUXFZCrCjH9F7lqF2GuIeGtcf9YwLw8qF+ndjFpPADK+
+sOJijRod5rNS2YbIiOobn4j2jFceQJWrAdh4M0agfS/7WZi1XtMjDUZHmzG7WcLI0GCrPIpwtK/
sSWhdcEY2JxZO3rdRyXyEco6p/g9qIxP5X/ruuvJpmnITzc9GNOKxe1lDp/8VuCFBdp1G2IyyY+D
vDib4RzsfOzLNvXwWZ1oNHeMkwVZUYa+PMvbqKxvJydC0DbBdtlJw0KrOvruzXL77eargBahDTfP
JX6f9h3ZqUDk3V5+pYotO7frI+e7ypfEienJ6+vI2v/bqGfwbjl8rG70EKhTUmvXXPW9cFvkmVJc
Z20I6Eyk/TlorF7HTbogYwAtMmzqbbRc8ZzL3rNjscW2M03DayRpe6gS4vHlIruyK5JpsnFQ012r
DZngVkRA0t4PSilixvB58dpA+zjLRXN5as0EN82VBjdXGyl36mixMK854DYuZuvBiIxsA5YamOkg
+x1MWlGQ669REVzO6UWGc58j/xt3UmZTPOo0LvsJvuG/rlB9L3GKKUBLOJwsk/F0xrbcT0hUdO+r
R4EvxTaA/wlAoRYkax7KPEZbwxGmPNEdEJV9IrMWPD2nQbWhRluVxCzqhcjPpCbNeE1Ngv1T26EV
C6FTFc7TpVlh0pP6/tDNDClp/tBXhO07Ue0CqCm9wlVZCcijo35CSF+B8m5P6zO+gZ/XjreNuw24
JgmEM3/27QkSRmtCQ+n8PhuuN+fHy9DBCCXdDUAdtQmjDL9wif0D5vxOyfK7RNYlxd0JELC5I1lh
LMX27ph15fz4zBpXLdovEfsw7hir0hUlvLJF53kegbH+T/ExwD0dwxsWBkZHAw9zZxVOJ+NWxFFJ
mxvzE3op0jXvm510k4Sp4N2imf/zGV1YN4T+jAEKf9i3eae5ESekzGorcN8nSVA4+0rycN0X6taY
4MzZ5TOqraBAANUOvRLJRpAY32Lq6ZhTFIcd+U566/b1WAVaa3VNaOS56/6HVlLy8zuuU8sFcIuf
MGYwUcwG7+RW08IZjWGvk/RXXjNPQ5hun/lsjP0ATD2M4E28KOcXkedX7emePNTUlGVlVR7zCv/0
4J5NEmhNVJkTDu+mqmHvDTYowoGkRWPWEsvPs0NI6bcCb8sE9zY6mFWm2AGUBXCY75sHj407OBNC
/Fh3q1t8l9vNHThjR0azkW2xzNWOvJ6SSIHPKquppYfkShrjjXuUac6vYWkNwkHoU19kSa3Ntado
xLpWwTS57ZWxUvHdQvbaPuVijOeczPz6DwkRu6pC3yr9tifKdZpknOQ1n5awzuZl5x5n4IDCEBiy
8NxeJJDs5gzB6eD7JVXIWbv8/8yyPDc0oLRgZp7mWFyLyCyiX51UshiJUbAfhcQcOKIsz1y+2O3B
GJrKjOE1CZSfIV8Gfj3JFVuWqmgsv6HSshYnJEAuPoAa91Cux4Ks79E/227ArIwPffbMOwYyci4Z
OuqPIRahYy1R2chJHRPDN9xgUI85VGp1XDQqiLKzVYJSl2X9S8eTdC2T6ZGywi2nVTTh9myKJ38+
jb0YK+r5PZ28SWbio1mn/V8pvnluJdBQmez1Db57/0B2TEOx0vI6yaQQX0SOebvZDCG7HQL35VyU
x5a6oUctr7KbOYOsgTdmeuFvq/+L65nOvVAn0k1fWbaxlGy7bN9yMmg6GQrk3QGnPgejyfZL7w3x
N+gedar9iyjomby7yK64P5VsMDGP16wl+B8gCR05pe3RR3qIDcWTGJpaZ7J1rpJ9MA52/XPLdpKD
Pbhvvsv1xzJJ1DD6rPqJqYFrH9lB8GpNcrbeCNuKi3QYzcwCNndl4vHcjvgNZUgq0qIALzz/aKj7
95utDDa1Ankk4Rwg5uc5zuqCoixXXsSKmtxI+hLHJNyt/PCKJ9kUGtCHdDopp+a4EMMjpAUfSnfH
XTQc2jZIk7sfAw7T5Nu46LHdFSNVh+jPC7bOd0gGtiaIwj81m/IE2IenEVpmICiiBG3/3cbdA4ps
3CGleF8IVNdezXL1a4PT3FWQ0+b0sV4WjBHBwvlaDOtY0oR9XSq2s8015eSDO9niUd9nMUt4SoT4
5fghKdnwSJNILoBEKP69MfjVV8jHzL0yMyxh4t2F00i22RVAx8c9ajZHo+9nW5yCtydqQqYOW9JV
UAsDgT5nHlTkrpVD0BcZBWf7c1IEtZCtk3ZoOIOwN0F2NkCJ6MlgNnAXR142vEeZMHyLnLBrJrB2
529gFDR0G46xf10u3Dp7ZyK1fUq50Vkj7fHQKO5m658M6+TTUuUOzCb/UFIALyoMMcYbDt1blGdb
HN+XUvEHW1UvwhaPfNqrO+muv/bsIAy5w6mzO7zC0drGKPhSfDn5Xbb91sAhEyQEMf5w4sX39wYf
biBosUSvBopCmlDUoK6SAxNGg2ER0UTXHkiCViYkqkvuu1E6x8csdbcpVZI/Ozqo4ouwkD7htrm9
hkmCQp/GxJg58cSzSI4drfRaRVFDW3uLapqzhV2W5gnut5jOQYebJ/ErQxFCkvCaV+CMkgKsvVsw
ppiefmu2XyvQvVfuwrk+7k8zPAyzAzL+U1D0zeGDuR71TJpkO57XII4/L5g8b04D7ikcKSBtsNH2
4QgSpxnuxoJXxNRSulpXzzrYbnGsj2yzo6WiYITfpVsi9oYWKPhGv0rWtYBbXfNfweuT0dSsz89z
R/EsCopSdmSK6BS6khLJSZXJd8pwLhfvpE3kLxjY3T/W9KMy6eRqCnVVtuCYHrmHh5j7GuTPe623
lAEyRdsfMs2IGRyCflth1s9QjvjFjrw65ynUMkcX74S4AZkMt8Tulh70as4BYQ0hTS2T1v3EZ2kb
ODgwMBR2M5C5WF6Qcpwps2V30E+EY5NHcMpUVe9//FrNcdBJdTlkjUd8hITAzbiY5bxNuqSmdW7J
uAtBKxes3W+zY88ep3tMIA+9oxKVjZYIlipLp2XILKWiTh2CAc6jLoVS3XieksDD5GQ7S3f8+MsP
YRYveN00gH3kN2XfOnqamow1jJoR23pgleGHD3NZ/D+YzILQ92CxuaQF5Yes//EOr48VcLrsZsmT
+BjxV3W7MD0fE+8mgUs5au3aMiqwQWtrEpqUwdwQyS1iAcQtV1MdRTjbN6WQpY5h5r6I+GYoY7F2
w/JiwBBniTlw0GwY7Afwdoa6KUkj3OxPoEmGeyazTcXfklz7q3Y7tPTNVPJVYkifl0NdY0Ofoec8
1rf0mpPz7SE4lL1MJuvuYvlkSpNjMiPQ6+vcv2vyPQdRWHuqNX3ux3eGPPAaGux6X9Ljeyv4qdAS
PBY3QjN4rgTlgP1luEBaPocdJaMaMFMJzgOh+NVeOcEY4QBzr0VNanymdlzi/hgABgHRiz2K/HyO
OToQ+9ZGMKbffSa4zVGdzyyETibbVBjtI2CoJw1ShfjWCjq6m2p45ognwfDVxlFF0IQM2/hiXUzs
mNCA/wTGRq7goZq0fVaBln3Twl0IoTY01uboKDLD70X4ivXB7FFwS8qulISHOPErRijlJzzIoWM3
4Co6dBAWYuiCX8sQyZMiL9iEjRyjzTd+07ZeIrH2RbaxLL3r7VEB5clke0+gRInkyBRRWKcCnqE9
TK7vQAu0rPSxZP8H9qKkSQhAlCtf8igfB5oUMoGhVeHtgklRKae1Vnm5dHVFT4n4oQ8/11cVPCDW
jHIPx8dEbz7gd8gpPqDv//ie1+TU9GHw3odIKCLoSip3GCIPT5qzQZ7v+H6A0eIY8fA/kNGLkyNY
lAeGUkY+6cQSZwubiVhj2or17ayaOjUpepovP/X5r8FIX1A6HOIy6H42BdJ3z14ONEbrCAhSjTO6
6QLBCFBma+p37x3vDuwn2N5mdnnYv8tSZpJQL5ifUrDbkjtvDCbYlpWfmgdlqcGrKjsFoxLmG55n
lS3NEuUyry8UEJUcjEFjtPWXJOUNxSQt3YOb0W6tGCrSNyri1ximcfoJHUWHfg2BESIfvT2qf7Lu
82nIqJpqIAhlyCT5Lqjw7j4makgIWKBe1Gp4jt5XyenQBhr1+mOwih3O7hd2ktZb7P1XVBok8oFX
2fEBixjo1a5gEyvxQd704GjznGsgZYVAdUvOMOU2aQaWVRohG2Iiw7XWeoK8xy6pp/rzUgOFmC0r
+H2wI8wFbhwETWW6pyPIVnEU8OP1/9CDE+YEYgBEhC6QsXJeQmi/Ufx1ZuoTKy0VfMxVn7R/QkFw
llzP5A1cyhY/Cyy+qMUUYyGvgdzFqBsMV2ObI3RZlUxhM2hwbCJRrsrdNzKcXlTUahzhJ5zjNF1m
l8KfSJ4iiF830OhEnoVOP7UgfluXJK6NsLqcTd0zo3jXRozNGWBleZmJRDY6myoThDXqO8gcFKCy
TLchrQUpFhtvDKUMH+gow21Kh7+4aL8zk/c/HBh3VbjXIXu8hlv6xqbRkRTKGRg8CECVGD3bNIAr
P6wNIt2gue9GTYGFL+sHL27npbHLfggGZtoMDXX4gWd18IXKdsEZDTrty3iQkhv4DIiOR6rN2C3w
4BuVsGUkAynyC/UKyC5UqKBoQNgFEorc4IqEfVbdO2bQtEQLkpJ/ZfzL9XydTsbxgsYOPMJg8Amx
3565HAqzgnvi6xzYwUfe3IPnWeEq9YauNS/GVZ0o8t7KxfLDxzz39aB2glx95v1bqcagIDXyHNCJ
qip1Ah/waUT+XG22ZjzyecCWtllajePzz7vGEca173khSKry7rid4Ih21/o+EAhCqAwc4DdOH9gi
PS6465EQk9wHRT52+XkZ+G1gD/eBIqGGanqw8cYd9S9X4sCmOxYLns4+xE0IYHwhm5QWbQsS4Ckh
z/n8OpcWHaxakwaOZwHwV248vFTq2MXb6ODALw0TyJwr/5RaCZN3+knHQlAzw9FRm5BAJOJGV/Ov
m42SoY2MeT/ehXzYgnfKo/nA++uJC8gF9Yn41sbhf0ETKi4eTOUYzPQ1pvuxTwgvx8N5inUf6ySR
xLsL7G0KJxLqlgWGA6fgzHrGRpefQXjVQV+EUenlRvc0dbbByBO6N8n5ADWs24xI/2gA9GP6h3lQ
D0GJ5KWV3wjJwD0UVFE47HB7gn25ggDHQr5bxDY+e5NzuOqkzMMsTldCmicNNyZp+9mmhHoinhyo
MqLuybtGkmKnogw7jsR8dhzlh47IGWS3+3otVggsCiqFC+WlC+GbJ9zSj2WfpoQBV9Ov3lAYiMNQ
v9tZbDanDDaiCnKf7njXO/UmLgUydv1aEuwr+yZf9QgLTDUXuke5hm1jnMtzLmejdf2iiBhLFtp9
cAYkEYgDuZrQxvOv8lSl2D73ac2VzVXPi8uGGYJ7zMfIXex7q408Lu2qEoIQc8J73QrGK/DmT46I
f3RTQtDCTQSddfEuWxS4fi2P7/bnJ3tQ3PEksfS61b0yk8Z3UW4DcUGvmS64+sVq93nLbBcOsXKw
FrAsTvMsvD5Qpkn8Tqfaz9iuMQLFg9dLn3koQVmrrNlPnbP5VsAwWxt+d4IyCO6uDwnq74SvPcwU
S+6ZqeA4NH0bKB9vbixXxz0N1kr8BXpJWqYVUCZnLEE19DHp+RZdfBwxPiMLBG9Lvb79LxgJe2bx
wK1OvWQKAIvTnGp29d6lPJhlbOIXRzI/9QdyDKkJ+h9QM1vLJJqjqYK3oSbK21E7qanBR1SnKX4e
LwaEY62Tq2IEoZe6l8PjzUmHEBQz1ggZ6TStHsWO7KI5ghS9BEtkXNJb61gQmgs6tj6Mc/5FOYPk
NEJstGJUtK2OA9HQdj2cxIgXBs0Kjyf858fc+JdiSOcLnnxv1rC3Oi+Ecse7SYK2NZqZ2V1thmna
h25a9IEJP0OsVtvcD5O0bpO9PMYm+evaUqGE6G5qS46gyo7RuBIh7/V02C+OrfVmzU8guRuA0Gei
O+VMZu55xLCT+QKL3/lzXoBsEgorcsTYMT49pk/QJ4UOKyjC2/zcKhtvBt6AYx9R5xnGe3C3nHIt
yS1DYbbmW9CKT/OzzjNBKHZSMR4VUW2H60qnTHrWnoYpEd2mw62Zd9w5vaZgSUAglL/dTT76c4vZ
sItXWq2g5QoZyeRva+eXDa8jInh3ttuRZvDZGQvLVQIYNL+gMEHuQtj4EHtRu3JkHwHjZlZmhntW
JqR2NL17AFh823yk0izXMy6r0OsayTx9FhIqukirzkIJnIH+m+n254xMDcSxnkIRj3SEPFag2r+C
J4homeWU/pf5hqpPoohOJeyjz9JS6c4rD6Z8ViaUZsE9sjA75pSFMavdAYWHjeKfqmtJHXk3ttt+
5IkQFSPVGopjY8+8vhwE5oJQMHnQpNlE6mlPBr7LIN7OKP8+2A1FjDqkqBMs4OjsfT0TcyTwK4Xz
980c3pqa1DZeZBz90ItmGSimY7yUWjy8TEhBL5jVR7rf43fY0XzN+1UVo2XeId+VG+LWwFdeBfqg
dPO2pkKoEolG4DxZyIwBqI3ga9ZSMylYhmeWs9igF/2bVlWZO2myRkXFhZS3BshtHY3vGO68WGws
xvoIheiDss7HJzravDTjWP5yN18RpNxYdR2FJvZvrwiO+k6hkqGrGzHC/izJbCRNktGXmU0W/KE6
SI65wmP9uK7O4JkQWesug5lLt48GPwCmoJtg3d8Adane22t2taBX+g7Shi/1s04w9eeALk1Aps02
ekAoU4wOoQpJoSzaKhIQcg3PdbiJfknj3si1r5i6gvvJIGh51NeTcpte6GCU1ae+ZoJ7vVvifp9Z
9irCAWRUF6BC7UygTqfqBKjfldDfA/gmKqFJpOBA75y2uhymOl6A+Q0RFSSLnBNbL/f4rskvDW1w
NA8teZNTRP9BGYRm9LJ2ouYzpVuM/Y63GpiWADFuwLnWxvhD+EtG+VpdW3XqSPcizdggcgIxBfED
5QazyMR4sAGvSi0tbuoN6t7teIy3arRHD45LPc4lmROmAkcMaouHgF6iuCjeahfWaACm4ZQxvWLE
oQfAcNYgdS9gbf5l1v6TRepZbcdPl5Cfu8HQXYqXib8BdK6JxtYTiTA3sTWXxWl07D9LKWS0iFLk
2vPnFxUcYU8euC9sI0DnNh5Q/3s/RkG/FPj37Ji+im4hzYYMbaSO819+ZOJzBoP5XPdynaXVknJl
duCljiUqvy0qfxg0nmwbwt8Ho26732Z5thyvYQRx1gWQxdEfl3+rcCKKLn2ARve3TuVBnz8HHMtE
3V5KIHrbnmn1bIhNrBJMLta3I6x3HGVGw6mVNpxYMkfvs2BgBdQu5I5Tzf+icuM8jQq8A948dwd3
lmH88Xyri777GCagNlev9nM5lA7f6uockJPYl9ZNTm1kMNtp+U1o7J42J/GFW74aGWFmqDqwdgSv
vO4DRWEy4i9ODLmwXTcVAlGEFcUyKBUwXUJBMjbIWwji8GHqmFfIu+dEmLvNxERfQ7uS98q56fZz
zjzZDiox0r4HbTwgzv4I+5iCCWPr2kptcI5jUM/cQQci9wkbDFp+Y31GqXGI9ifR7j+bk6X9BDo2
CEFm+dqWEXZ0i6RGzDPlFq7eBBAJAVTpkRpX7Fw5BARXLpmYOPAu9fHHcOY2J+O62pQEj4HfuoN/
Wj7LnxtM7Ksdun2veJHfXkt8/3A22KnJUlqIgXUf8r+uRb1n3urGVqleY5Ex9GVJjaE8SLik9pAi
rvPvYrt7PUgKIZAquBYxf0uBwl8gzY23n5xJ5CcXfPBWHrlhzbCL4JCJ8+Gdt+KOMo8oUoXO0KLg
YodO64MJMUbDNAR4LJJ/3/yPeRegvxuKyo6yKNc1BvvP7yLm7BbhL4hZfz+QYPrhZ5tNBAJP1FuA
kWa3IRu9WwvEnPNe6MSWdjZsEQH1N4o3mvJ5+sNl/cJBWXHcOVQtfp2UVjPjvj/cj3zG5e0mdXEp
TGk/9OfdVh56CMkYNDn9wB79JoX+zuXm8qJahJUkrMXatSbe0oh3ojswScX5WzU45DqQgZaoR4hP
7rEDUlEU3KaLFL911CTr1Cm46Q6H0aErIHj7tXMMepCRCgPD7DUbxNehqv2/NzKnVV8wlpQ63OeJ
8CEt0FX6rdcb95AoWjJhKBfW2ZEnOUfqu+5RWLS+2WvnhYwM9LSXkOFEl+9/ihyzl/8RECyvL+ad
I2Vc1/aKH6E1DaSVRBacE9fDjKbQdVdyABcavE9yLsgMPtpqMOgbxKQYQljkss6JgUu3OGu2Ju3d
mp+sflgwq+SEHRvI6J/0ypYB5ujPrCLpr8ZHwFRh43NaLjC9mSz7P1hVfMm0mB58viKxsmN5FCRg
7cxKXcWWoJbtVJx+cO7I2DimO11fLNdoZtyZ8+osz1oyXpuolrOCw5WT6tl9qFaZfEaSUr8W4Xm1
pVBi67qPjnl6/5oO0AUNAD6luPPlLiiqHYD/kMfIBURCdCt15IrEi+pIDikx2b4BRZGR5fk6+YLi
poBLsorM2mj0UfVQ+ZDzFfk97B2GpF4uTVeF96+6SluuziU+7LhWtsEk4efQKVT5LKN1eIAZa+Ny
Tr2Zw1lYJJL45obDl3iO6YB2Fr27gmj4T39Y4OcCIy/aNF8FGBDXenTRYV9sA9jsDhkxzwuAudSP
63jWvvHIhCtTDwjPvyK8i1Jq4b7M1awh4WVrkmLT0Gz1srAhMlolKR22d943FdCzlnY43CSRbVd8
KOz6yURE2PchORzu4yRR0KodwZVJlH2TLoVWyiXWv94m+HCBTaZNVD80vxGqEXqPN6/CzHXvp12H
8GPpTExNAgNJONDfXETr36TDjSu7K5c46Ch0UWJI/7lQ3mBrD5lFjtBeUEAjdgbuV95NvXm3jaKR
qH1SOjzEDgcvNbFcrFjqlJSaqRyhrbFR+tkpPFTiPr0Zk37AavVWoCP7BaWh2uNcwP4A+BHTbU4t
JFoa3n3hUDbk8+M5sVgF3NDewICvTAYg269ksjW5mS5KdpLRDTHerhcLrrPwEf3Qd/QNItOOxY0M
WwuorOfGTxW9WC0jgK4ERb8eqyACQ1BMJUFzBpoRITkoVEOjWwj1AnZvlQEo0VYAcXLPU/BWyqLD
oAX7o0RA4vwrd25gPjddFDxxR4dn/qh4FU1HUM9bYI+Q7RltC0VwQJic2icF3D0+IYLpc13J7QcM
LV/2SNeeKP1QJcCJVGfx5eo3hJJOzfdVsmjrmcsLxXRq5EDeCZgDv3WNRZUqXKSlGQZfL2CpNj35
IImXbOUdUzVjSTAiSstu9dF5E/Srv/T8Atjy8sahks0msgrD/VeE2eobcS/sM85e3ccS/nI2mTYq
Uy0nCngCN0ePFd01Rcf28TzGfUMSSTSK0OOInxV2QHH1TGbP7zsjPCYAY1AMMNWdL/QwbG1fApY+
ttK9q7UdvhuPyoKjHr1cdYK7wnS6LVAkjwdLLe1Cp/TizE/GnTgFMlzr/LmCHKPg7CpN2N7wiawh
deBdYNpXVexRVZxbwESX43msY6bmPT2mfb8++rTKyJpU2MtVheFRHfmT8YoVqw4cZUh6/ECDyWYa
OiXJqlIXK1s5/HI6r1IC2/bv/X/KAtiOBOWTzBu//TUUHCS0PC9oWOiHovlpZS+J49Btf1lo02GL
ZAiSHo0a0vvcmwG1FapAbfEiLT3Vx9630zKcRkOZ1TmvBqOPoEUSzIOyxUdqSK96BF5LotWsKu9L
SxiYC1+XI7Xxoop3Dom55TRcLV2kCAjPuDOTB3Rm5wtI9+MWkCZwFF+NB2/RM1/MM9OCHK9ZEMCp
yMZF3QDNCXNjurXMxlo56eteHCKMN+ojyMzifuK6+/9zYyIFglpKZR8fs6YFosvXno4U9UfKNmE/
lhHPTBEZzcuP61Z5PO5vQf/iPvhfekaEDBROf6yE2Lvmu/MFauJXxJOQvCVsOTMerJlrwmfbBk6l
MJNW1svdgUi2lD0KOR01/pCRMIS1uEQgdNJgwHPsmlXA9lZAt2gQG+wOR0DXZK3SMC5C+/PESM1A
BP442UgwYqV8PEenxx8q/XxLliHDKm8C2iN0YdlY8xBvzHml7hDvZYiDzBR8pN19enpQIjn9B99B
vreHupbbcVekswtM2Iq/++ErwnpzHkWztLKskU+adk67GXmE0i55qbNtDOz+3/7D5HIXqK0R6g9d
Y+8c1yqazqDmqb0yDuPSLEFWotR2/IxB6j2bdY/971DYsB6PJmgm69E8mxigo//+z8UgGTpzWtYL
avAy3LiuLiDs5WXjCC6khFWv5E53iM1Mf9Ck5xtmKMsFuZAW7aLd3Yb7QMNPx2eYDORkHnNFiKcg
l4f6x/ie7KZugsfgsApXnJPryiD6yuznBupnXYNRJq5kGMSjs8ejv6xaqZ+aVvvr78QZqJg0xQjN
rsRSY76h6ci1dezXn2blDQHD1sKD9vgDiRpsPWvY8d3XT80Ijc+4CwNAnYKJNlj/LX3lnIlHwU9A
kxFUI9qDirwI9xYafAtVyqxZFx3i2n1cV2OTrc2tMx+PFYiqsIZ2H8PosTA2E1N1dEA8tCgzGXOq
mU4mAdl3V/3zcQAOG1OAPHwFAqgIlpI5ALNvz/5J4s4E/QMy2eReNmBGf7I6k3GgzP9SmLzNV1Bs
V6vWvuFTx4o3qjZI9N0mqfYh+pwBNrLipgoYCyVGwmaWlJvq8KCADmx5CgzxQKXkFKIyy4TM4/EF
SBA+Pg1nHSfruWKMUlIlL6gfAiPTPsuY5SD94fVAdxPExTF9lDsBtXRL9Fxkot95yhdpAv9ycUiQ
ZiuH0qGcnuFSF8fJkYf0xdwjkxCDAL144wGWk6073c0XbyJs4GquY137142o9hHqg51EVgSKeJhE
OjRaW8S36n2RCHS4/j//GGaOD8i/avRHYlkNzkEkrDeYzMe+vTeUchVf5P2nm/TBfzD4SlLgkZmK
ppPyvqvOwW23iZZyk9V7HuXOC9tcmfVplpTsDA70djRUgh1K0WulB5BfBJnfIGg1egCy3uimMjSt
pBQHfGk5kPLVR+SietLlP8QyhBrHpiLyRyirKrd1g+FD0nLJ1rZbMB9k39mE3lrTBwugZYPwjGsQ
gc/CypiDq8DGRkW51Hy1Lapt1AUfWTd2kIZ7xAiXEoRr0CIsX0046dThezGK45aKPxMOOLU3nLZR
Yb1lDJZIqca0hqXDg9bbhd/yStIV0VInRnQyotRoxwhCWPSBq013gFbneKR+JWlFLrqpm36LBKVi
f49tPLQFPkwSx2y+opegykt+g/KplbsM5g/bWcoiv7Em6Bm6OjTLlNwKHCbIMl71S5j4W+29DwyY
2r2x4cw7MQMjsOulV4O8aw6QFoorEdp24XVKqAsp5UcLSw597z3nEmvZvGX3FLgU8kJmbFUcCUv9
gqOhtc0FwlNUT4jrmrRiIck1yslCgLYuDHGcuP8M+az25CBtO/uu9Y5O5OpDfN46M9oAGElD7kkZ
4T98tadlt7nEyf7ZRTEVGDncUi1+Bse44zTYnqUBer7qXgTh6u9b+nQiAbppsSTXm4UygYAe8AM/
QYM0SQ5kSgBsvmCYcDH+s9v+kZWb8V8qnVqJ6J4/1GcMuyQG1lyyJEhjXG5KovtEePvrh/3xkjss
AgI5Xir4ie5M9+C78FziYZP2SnvUlnX9y1IByIH7qgRSWfQ7zSFXrGydMPq1a7D+O3VzhUJNuzpQ
rUh6GFWpulRsHsXwBw+WkemVIs9D6VC+o81Xs9a2d0fpzYFIxUiQoSZgMjqiSwxefT/wbD45vDPy
PSnxUnoT4M67pK/36thVMf7X/3iBut5wuaNl+ikYRvEJFNYpgdoVWVqG9BavlTsUCpa4zxX+3CJ/
6h/nT/LNCan6pEtN+I7iHjpeXpDmO1qePKg8SyBN5d7ap8EpcFXDfVVlAoLmn4psvW5UVXVRw+4t
/2YG2F88llUypU27uvtdvlJ/AAAXJvReXD7A8znH9KY0Z6DKbIGfN/wfRa+YN0UU4tAeLOeFMw44
CZBenSitzltGsAjBU3r7W2Jdid6fda4KcYLwTEU00SraVmzDd0MnXfUHyOPINyo1XYyNBDqJroHW
aSH0dfR1gQ+rqmubV8CcHC4U/P2t5LY9XiLPdoXlvrNnaECZ6sVGoUKSbzKjk0IA6go+OhIVsMr+
iOKejSOtvbHc1XdsaY2j+7A8mi3U5k/BjOA5yj9zoJQ48CmsdMM4FCYRaKDOl8+/xuoVQhvRVw03
22WSNC2l+Ljmh9E3Acj0wMZaLvdyjLW4PscH99wriGi32FWyJgODkGvUMi8KVyyzrut5BFtZes21
MT+hnu/7fvAK/oZDy7JWhH6I2JoA7UdEFKzFU1vIirAfPr1X3+YDH5KKomxWOvVo3/3suEvyXUwh
ANvz8uxyLQIc6COQPcEr1rCNMTNjyCf9KZJ1FMazC9Ou+PGjwaO0De69EuX9rG0+yzeZDtVUSL3j
nvxDN+LWd2/yD5IqFMajCGCqon+M1gg5rg9+e24v5gNjTVF+GPLSJ6tvTIdua9K77tIKqlBlg3aq
7rxVIu1Y2dhxQyE/JncdDW27jJSx8vXVMeKBJ/NA4aX+j6f0mLI9xxrUBhXK3RVsfe8ClwNKBUl/
VbnzH/d1wQS7p5WpQhdOSW/JQ/eu5kNQo0dfosz9rStP4IsfZjTDou2DIdnF8n7Ee9GlOMz0S5wW
6nhHRlC4iIJHqD9IiBFYJXirtzyPdJKij+544v8Bt7wXL9ClP542dsROvzeQJ8drIe/bHLo1AQxl
hWe/2AW3JmQAJ7slyOqqCKK+jail4xPEHG+Hsn5GczEAqmGGRJ7dCp+qJFZhLKsjQpbODAPWHSSG
fCYBncOfHlIDVW+xS00hM7OvPxyXQfa+51JvWpZXjoz9kAIY9D+hhiY+QBvKdEuRiWLeGSlI7ljq
9vnbkcYLzQfIHymlTtLsuCjg3UXtEiiH6MTsgmle7QmjMIGoN5uKJcje7Y10mmMwkQr6A82+nD9N
3uuV1EbVl0SfuBLy3amhPqp08ucmF/uJQSFFRuE7qlG3qqXGb3ovyEifukMnf7S8KMWeDNLlxObG
+jpNje9ZoXJFXKn8auSYvBYqeKJmKyFIU1CI/ecETaAXlPC8YwaKxUDXnyFhz4Cedfd4nSZk5gAs
w46AeRW+Cdd4EuI2ioahikB1+K+L36Q/lmI3R9R67TqXKweJno+zZV8S9YA8vDtJTutrXJ9CIY3V
gra729RzsIua8YB6oPHEhyUkLlvFBgFbxK7ZDVSC6RUtPt0Ej3j9wteFfR0X8IvDaRM2Z+iXqW1f
xNeHT9SUWQ7w2Edy21+hszLNJdNDyOCveV1tDSdD3E4LqxA0NxEeg2Wby3wyLXp8GmXT37Ed6ZkT
yt+GH7i12sxiD5yg6G2ycbbxxqedIfQmFq/ScgaL1RDoIHHbD5MJ9l9fAuEuced3I2iSrbp7wOyd
cdPTw73wtzZl40FQD72JwV7ienhc/P4H9ctypqEwM4igXq3c89qpUMlZFAY/GI3uS+42QeEcrHUy
kw31coR1B2TnFDCAC/4x54DC3JnyBLJqxWovBfMTlA7I+U7Z3JN1nVVj16Re4ZMLXdCDWYB6Dlsi
pETVC8g1UAT+T9hPkY8A7JCGnGhXBwxc3/1B/mShQleJhPLkxzgONzLnfh+nc3JT5qeRaHMy6eTm
ZoMyF9VP7LEOFrcjNmW5ny0F5X5k1xIYfvEoaU0yxM7MaAJzMvOMyGVlNHas0fmDxdvEDjpx7jv2
c6vY6aofN6/FcTZFJLAJxuOk4RWETV2kPW7PQj+pDl72UZDz/PAbP0SKVsKLck7k5kdsOCalJacA
gHcn81gWIG3EsI+AnpjPP3TDwY1Lv83/D7AdcYQLOLdnZrMGH1yxQRdKXVBSbBGHy/zTQSsS/8Xa
5GHLA+2odqrkBoR/z6ernEt98khXoL+Gx+6Fws+sERTIg4eFuanT0tgfmx5SCIwjCMxjpFIOxVOf
myS4p9tDHwwyfnJZA0XEMZfDKW6GEaihXII0AQqu/nDL+kLHvi7hmfmygenUQ5297fKSGJCztvgF
fYOjQt2GO3i0VC+cpjWXxrfUJ8pVZvfnIX0tHHeRhgHkm1w1Kk83ONNLcw3XAfURiAckYx/4IDPE
SiqZuvggly6SZWyTow+QJq+76hdZgNlmrd2KyNuW/z530NGm0f9WHaVKLoUsECXQd711D2vBPRxq
Si3TScAoWzEcngkljSiZ4fNsUY9oMNq13zH4DmKFSK5wdMyLRJrjX0TYA2FOwa/B1hWs01+gDA9S
QekZga9wbmOf10JCHS6XcJCynMS1aCTg5vIFQnr/r83Z/pgWcQ++8A91Gjw4lu+cUGEzV7A96fdQ
/XiJTjLLm4qJ+e5QEGxORXc/hnZgTdNKtQ8q/pRkrspCs65+hhNvM2GpnnCu/zjUkbzxr4TAiczE
M0gVMtplS2Gb8fMW5xNhl4KvmnujNOQ4hFQxczRoURMHiWC0ItrRxDVvLV5RuO9q2UhCSpxPVY4x
EmQnweKYDJuoYDgLrPNjA55HyjRRkJdWux+e5YsYsJ10iE1A5oI5TSphcnv7u/bSh9K2dyme4H7t
NCD0OuPIk2vtNktgJ5qeqBxCN3y6cS44bN9rOdEODLrgKulgC0PEnJrsFPUFINYmqZaT9dwLQhP5
qv2DyBCvinpo9sW+SCXWrLWQ4jLNUoaoddEiTXOLi66Anfx7xrCPhTomOYo43XVEod/cgSrKO3RP
Ddt4GtlSS77IwY9CB/LjiVLPMbxizayR6jcZZa+Qlxq1gnXPwYRFqpS83C7tohEdNas0d1GCXQDA
Qc+QKt/xWDQenG7fkYgS3SGGc+TeFVo5j6bgx5RECXRTJpRgBkmpHFIKSqmi/k6JjUm+XKG9dlB0
KAvojZXwR1ZwwrqOoIMNuQqjzhLjOrMosKyxhJ4TjviXmqFzoiS1jmE9/32Re2ZWoCKlpKjZ2iKY
LCwT9sTKmqQYKK69OrWe9NVIa65lKd6DQquyjwhjZHMl6Mg9/dgjwDzXvcOW5jbmDNlf5zyAdKEz
mcls+4F2B9BRvpp7YJEHOv4Ne7fyy8Q0qaEX7LpDkjnEAa0+9pqfsAPVq+2KBERA3I71P+tc9I9C
1pVvX0elYQY0M5qKkF45Tfz6qHaGPBa83DblQ1ZvxHOh8T7J7UEFjxnogXThdBjU/l4bnNwqr1GE
uiBwUuyPeQQ15gq0rTlJ9jBxy04POlE+hnE19VgZx0X6RrBnvQVR7kU7ID6wPcuXQZbqNdCyayq9
vdbJwjJEg4TrPdBefKbYGFbg5DdQ6Ps78/OuVcne12D2fhCc2xkUXWxoLge0q9SELqkpGoS8Kd8f
TLIJWVOUP5ytaNiwV8MeIF5luz1gzbIbSlhVJW/IpQ8luXzlwe1G+1vHkZM3pix7r88E+tUu54Uv
oXckRtcb1KL3G7xKfep1NPZE2x4OJPptLWBXerk6lH7VtLkXTsRKRMlEBf6gmowJzMuJW34DTO0+
nd/VOd8QxOr5pyIOLz97kZXne+08aqoxGM+4YmlKwm38Nm5/oyKlFdVQ9EBfxxQIBHOvpt41H2/q
36Sh6UrsHO+W9VZdqmtJunei1CgC9/MO59ESqZk2X6i552A6njZdrpMdT78BTF6QMVSlBqq7Js2m
SnSh3EMD7r2P72wfdih11gVt8PQVnegJsA+ju74kD7hhNiW5ENqlGKdkoCT2k+PDoOSu87QbMEWr
bCObIdugvaJR6CPLorHGr7HAV+xAONV6qAMYY0/yB7AIfxlwAldqPiGPg2JnPIOD3Ql41g66DBx8
jz8sW7x5MP+qmSbv+Rf1WT8WuKOqw3puZhW7BjqsjHfWoS1pv8dxIefQ8xjd+9ryyhC6iOGXqCAX
oBAsD/1U2UHC3y/spErm9nGXpBm6QMB5e8ygotrDVZRWSyW+0E+sdWreRQO5PJ/odO2Yn0+qtGC7
w8y6GkNDmaPVOraMLGyUPgM1GgGkY4tnTmBXQKxoX0UCop2pHzQr2SRFP/ClUqMuR4VV3LDhL2ZJ
hufwtQ2owhu8smORoDnZUNc0zJnAhIn2lb4gePECtURTpJHk7LdPXIY+vUFiudEb8WcHxoVxgZfv
RdjxJbp0+Ls1ToRbzApXyvjsSbiBFQdSyZKrx+4nSLcT35AeKRRdpWJ8GzovlugkaT/EinEyCj5z
xOuOnQmpqtYDYy6SgGyBd2xP/K7QrE1yi/fpZ144Vu8pB75OA44oCnmDFRpgrUUkoer1IHXuohkp
cVjRkbZQ2GP1X4h7wypJC6l7x7lQEwnlrwVN3XokdzfWxHFT5P67Ol+l+0PqcQQDVIhewQCkvLWl
LSDlGvJJfQR8LHeCwpxtI5iaYTSOqv9KduO4SviJvNzriS2J15rSzPn3RyNx/KVISTXwHqK2Sjo5
jwNwBvB4HIBFc+a7Kza7JG2xFNxHqs6VgIAHZ57eWfSI8IStaNlYpvbcU1euiLGy6ir+rl7AYhXF
CBgKLhyElQoGyqT/ag6ASnJqaXRmQpjF8W+0PJraDidQFZP71VHMoq4IhpdDV9U4AdePDaCOWVrG
vPM/VfdWF7S86eKk/9qUfSjsg9FA0SLiwsLVxnXvbAbzWAvjzKCJ/KqP9HgLBhHGp9cajykiCE3Y
k8RbfL1zoZK8VmJArZSD6WcE2bGmZ1hJ9wK64rsSMEOWvumKT+Z8y5ibf+oDE3ZqTacNCZJKsj/g
CuilInw+bDeIZ9at0tISfvdFknbBqvt1ckw4VtU41VFL1vcFYWbb/K43L98r5nzXtdzeuC1IneAF
x5LhJCwluaM71qxlMkXN3j1zO2GBLb6r4ugPPY5WszHUjSBwhvLKtoXo+ctaZvlq2keKoLgcu4l3
IzXoDM6oHt8Dob9XVoM+DTULIf11VPvdCt2wjejPKZYSNHeGIl11fCVPjsC9fP8Q6cNpG0kZq1MO
vbME9k/KocYEiE+pzIO+9YasVu/MO08wR5KU2NINFrpWJkAs7HxMGfd9+72cbPHr0xocMkaX105I
GoYmhNDuFZQmVOO3kIcL4hkX2b2J2AkJeFNBYOtDG0aqoDahKRKY4e2iR2iKmwEid9QzDO5pYXq7
Ae5EGbyCbzuDqLN3/cY9Y46napWVjhQKuj8Mp7QwDHCqdZm0XJ5XqDqZm+a3UAqbCgLiJ9pM9pqE
fI5lVJ7/OWVuVFTD6pkDqq/ItBre+VsSP/UIr0Nhd6XBTO7YePoshZOaiU/plnaN/skK1YT+jNXg
/D7zDsO4benfeqjHUh1ABlggRWmKItPGEOGubMsPljc9PsMtpwW2dx7PavElfHHKjgViYO9NkNfG
xsuHwEvpb+qw3jZbHzSiHbN/U3LyQGFOlAWyn1K50dqgp5fyxWmZJVIicVRwdsfk/wN3hS1yXiuq
JoEv+NvZDW942ctOt9EvpDUaV0hWAwJeoka/4u2WzxBd8cBi/SLzsJQ3rAdKdq2dh36J973sRkb8
k8d2ezhEBbFBh4OonYYmFL9KiWsQIMw/iDCMM1Zv6MbIxy3NgYKaX/1vrBcNiILRc+FBaqOgsePG
S3w3gn/cCLrFqMevgpsKsnyT4L4pG9DscF6XOi/cLCaf4cJY6imtkyQZlQeXKwfkej6KWSVFBLkC
bHm5RueZyR3zS4eGM/ZTqT5GtIRZ0nbv+F5LAZw5YoC/K08U5kKHlhHUMdnRbh2QcicCdnjN2oCr
vPK0Z4qZG+AVsc7X/MbPuwrXLbsYb9vox52XoZvcQDQl3yb7Hx93J/Qtj4mld91fnqzJmAXIKr0j
Q9+qmyz4diNyaqYuK58agA22KTE5bzwIZyvzq7y6/Sw5ZYW3K1mvX6Upd40U/fFfO/RygYJPvbgT
e4M98Ap0lqq7u/i3htxIRpTODblZkP3nBZ3Un6ULQOPTOYXqsx08DWcbFspNS5fLgcQNLwvAP28b
OSh7lWpMdFhCLjUDGGLmcNj66vGkvy0f6gbqLCvEAUuhsxKn8CII8hjPKm2nMH/yzTT4Y/an3MfF
Wv8/QFBGIMaEksGURte5qTqLk9aF9mDI98Ck+y260DbXxxD6rW7OEYTGQ63ApDdJ6Dv8avrQnVqs
xomXF6aePvwrzZt6mDV5zf29UU+aFKDMFDeATQ8F7OdmbiImJ0TZqV553NbQO0nduLJkpAsumSdN
6JxHj5WwrYtOQBWLpE8Gx5l1Z10THE/6x4PJ1H1DGcgu96m50WFWXNXwiZTjaGb+oVwztlV79rkZ
0eDl5zg+6z0sWcU6JshslvvO5zweKyPgbbH5yicOGVwrwaSB2wV73p1PhqGY/6/Yojy4CdsncqTh
Bh8bcdHeqEZq3A47Mnch7d8BK8n0pbjEkH/KLDL9xdhFFulnCUSV5E7MZTMe7D8t3lUuEmJRbqP7
pxziF02nkqyLwp53IQ4xHWajTihLMfnmtymIulJDTT1rL+f5l/H07Wyvf1WTHnWl+Ll9S2uZJb88
eqxx9piAOXjiYrNm9uCs4s5SNAZe05NA5S20klwMI/TPCeETwrPLAs5ILmk1ui2p5ZXoJpwKCCK7
YYGwShJ38o+6R7KVXi5BYCFuUkCDYq1fglosCEoNnxbGcoynytaofpqnuT3u0ZrL7pmj+XQ7QzLm
k7ZTKM1sUqxYWOhwqdKWhfhCYq7DEDJsdryTZ9xsUBwNWLWnSysO7VV13tFfQy7kESUXfzJCg8MS
X0WxkFr92LkIb0I03wgTMbmXKUfOiTPAepjGcAgYGHgucWqloOi4USfaKJskc2z3ekQK4yzjDpTb
/s9H1qx7SaB0PvVOT7VJhP2O3D9t/Q2mqGRXpVYG8hQlZgCksYeoWijWb4FfuW23d9I3hUz362x/
oOOKO57+LdiCbWAYwWt1LMpbAmUuzZh67ywsKqMIskPiHGMOy7ANxqfhsRBdTKY/LsLUmNJ+4YiY
fwc+Eof5Xh6ij7Dyu6FmTuPd6IH0yKMdM0c6N6jyLAmgj7UqIyg57kiNv0ZR32jqiUpk6inpfWjY
Wnj1/74gAZG0PQMq4xnBGnFAmupPIwOXxs6av+UuNIjS6c5DYwe1BQD9AjYgbq+1OKf3ODn9Ff/N
nbURuAJGetMJ6ObM6OGrqSHcs2hrbZnAQTpuWnFTO2DwozgAbNscBwFMQeZTHkJN1Y3CfeuxKAKu
XMxx4TNMehS3+0bbRhLJ+CKI69raCOuqD7GZku0+XzkpGuqjODUAek+i6kdiWPRw3NRweTgYRudd
WbGyqwnvUIikLcqEXoOo6wv0w6NBUhSLOgTpURfGq+j4ENgG3fps36/26GjPzV8UClTW+uPka6Cq
etPnlFhQOLvVgeQ8Brney+t12O0Yr9syCnEVmDa6z8nDbr06bS8cp6hM/cm8AN0ylPeb7qDLhr4A
e9AHyUz7QGqvJMYBDOMDc4Ns4PPNPHK0ofGmfdLPSvW3lLlJUTcwLXUuZNpjC+ni8XpSzfjazXVm
jTkLSl6Oj+nH8n+wHgZCOhJgSfZ3Na2W+NQf1RYP/wSzP1YSxV+L+gDwbc3XHu5yysd8eRQX68Ea
eK73F+R7rF6AHy9+Szau5+Aprngr9CkA64uFghgyzv2DWO+RAot4wdYGvY/m91Pm8dGAk4WQTZ79
4zIKRvIT/xjgYHxCswkmI9Y758cXJ8+wghsEfWRH4lD3YjbF8WW7yK4Sdf1KVKuECURY0AnpuDw6
jgmeGnjlIOCSY+UL96P3cBIf0gZMZgt0GMS6QvHCUMqgvhStaPPAa+yoQ7ZCGXslf7Jso8Ryc2ll
6TCp6ZKTar7HxoFz1eHdbyLghoWM9CQ4bCzCDxsfdgWBWfwb0wUJ/tljO5gO0S8TzBlC4Zkub6tR
3n2jeSedLNnrFe1xJvUDFoWeJEihZHws9n9q2TiU7JIyfZe7cHV5lKpbQGPVkFdy7V+tf3j4C0Dj
54IyFFd8lVsX9HwCniEkakLacIb9q6b9pFnVQFeReGtxbrzKLdseyqCEDPjkgHPhVoDlx5shn+pc
e0Fb2QlERbg/kgwXVpZEQsakfLQKnXNicl7gpwHGdJffR1q0XLt2GHyGOCivyjbpS/AfvYKZV5Nf
V/I94/NlfsZZT9yyrzX5s/WnjqFuXSWUilivAJ1yE1Onc1K8srlJkcC69E6lMCROXIA48SGaTH9G
svd0fd+7hl31Px2Wx1G/Bc+zn01rWFLv62MKPHAXQ0cJs3dUAMcFzwka9bNtQ1H4XNnSsEYsbOWu
0gs3BSt07EeDC9G8OoknLItEi9k1X+D7UVdGjPIjPgQkFbto3xZk+d7AeMsFuEkRvF+C5AyRITKE
EQMg5DQng+qgen9lRrP+PNbOrJZpns3oeYgY0iHDvX3W/nGVWCB5s43wfbBTDDnSfM5FVetroZO+
idl+rMY5NYS7iLYuCIp/XiOj1e3Z0yPL2ZGtZTpGGlTN4RLez04MpMFAq3lhQhwLpm4vXJhQS/GI
Q8SmVbvgRWi/cTjVeAzNrNRQeV9i32lRgbQ0/Sa7jvZo2yAWEVirrEU461A+joSZuIh48R44rHFX
CG4uG5XAkxIir+9KDDM99Jzs3qc74qO0rNMvm1B2nhQjelOmK9Czzo5gV3+4vV6f2GYWYRwAcw1l
F5ENcbmiss8WyEwFLAnrAH8cmI+mKUpIR/UhiYn7D86p7u2gHAFgSp3WviO+S/qtwrSOAQc/HBnx
NviZpmB/1Ylspp1Qc4WmSa6tCQ7XCMyf6QIvse785QCun61Q3DdgASMPtWLhNt5y6ylaDrt6R5Qs
2n9w98Tgh6NTxgvIR+3gcSqMHc3hJ+3I27rfJsr/wbMSmX79RglCHuMmLZH2y9OmYcdLLQm8vX0N
pwXiAWaeQJdohyxIFnSIj1fF3qW3HbIkZftKIZMDWDeaOwKmiEPj7YL2KUB2WcvwQXFySX0bFaMU
0WlMX8pxvHQ9/aqyenh/l68pB+bQwNYzrpALo9lfzwiHgYL0CWuzNaeXa+zB+QH4SSIrEmi1Qctn
US89nt9lgNArTWMyyLFld09BaGklT06dH/Pu8MuB/8v+pN0WalGC+vNA61QJSeGYGmAlrtPMEy4u
xmMO+G4E5Ibv9ti+HlKXwiwBY/IiIdos1OlxK0ZPiqE6oMUzIAR8X44rZgg1yiM1u08+uw0D8MOM
/dbxvmUvYuLpF11yG73WOZp+csePSnKYhzwmRH5l+M59uS3C8hjh45t3F3+nTOxSbb084rEoWHIz
UQzRu6hab35h04YK44ELbtGeY68AMZ/MREpqi6PuJeuDS4PLXxl4r9S5HKenBUYx7QeK1VXlmDe+
dNYhtlOXqU5dhkC2JuiVS/3qJiIrehzmTGePpRV1kRxVDtKumzJ+0RS6hpA/ian7S2TxnLUGB00G
vPcP2yU1sFaZm1VVGUIxEi3OorkdmoFDeGVWhO+q1AfCn7mwNoPkHxLa4TOE1p4orBq271/5uhU1
4HzL0s4f1raduIvaEedkpZVkBc2t51kaLiAE8P0HkcUcnQp3EKbVqN9y5aqkXvjUI3UQj5N1Ca//
xfn+8axHao+LKDqYjHeWMOaq6I7AgN8T2Cs5ebKmf+I4PqpfZuPRHrV5cTCSZDlCnCAhPPGEI4NR
6Lzw7bOtQUOdpFPoGcJGAGJnGADWiGRaiDSBiD3qnigi632TQINasdhl86Wsdg7gqXZ6OOUcaRam
XrcNT+IVa0o2vUfpnkFYPnp2KB20e0TApIz90kR1Gu8Gm694HT8UAdeIXyYx98uEDnHTPoNBZwLj
o6iTEjvWOIKRmQrn67voZUfdDhHqPtjUFhoy3IXmbebfJqNcthUroKTgRPEZJ9dLVq3mpFLg7yJM
+LsMPH3TiGq7BEi5D7CEwVi8wUMLNUMpmtjxevTE6Jnqxr+2p3NFDE8WstSeJHQN/5fFep1dioP8
UQbpMHCSWk6qQ5plw8p6Hv+mj8n1F3jjzLxQOo9cY8OKti22lVbV1AP8Coeak37KfiLfqk4RSTCN
7ag8RBD5qFoq5cQqgDn3nvak0Gqcr3BWmDzbUwsiMRjEr6h3F3+t9wiLhelJLEomEPDL3J1ZOU/b
IWCdGXzhunGVAZOLoBA+VtyjU3sDkF8a9Sz++tc0qlff9ZXZNcqCIeNg/sHNQQh0IdKRPZ3vy/xy
uJoGZSMWZ3BeEOn/scjm1lUx4i+12mY575Z6Kkzmcn718jzfHNTP9czvzbKgkEpg7V5KJw1Ujrcb
+pKHq0s3j2uN8CgFfvAN2hKMkJxePKPQPxxTuiBqh+BWCIGWCJWDEwkdU0P6qyK8z0AweqbwPnRA
qxZFNYk3iauSTwtnJwEw3LXY4GGKMNRccu6Kv2EjwlUPxxbsBs3iUrL+KkImwliCmFL+4/kFBSE6
hySNGAi//MIkKqo1MeuJOg9TlxWQTgg4rmNX7M7um9RhejHc5uENOjWVWH1XPQZLR+CCpBm8570B
4et4o5COSDUKHJdKFUk4RaD6ZrG6Rsa8l4xHksTkwNmKMgGLpz2YreZoKNbd9dT9XXb9guRwAas+
Ko5vHXpLgBH4vgazKTgFT9BpwPKF7K+7EZM+S2RJBP/gcyHyIWb9nm0m5gycfH4J4lPscncRnjrZ
3zpPQTcjMjmE/kubwyWu8jcubbgcehoqUpZXvayKlAU0Fc/ru2r8pTY7Vk2S2vclyPb4s41zDpvz
JueXLc6yal51IKxtiVnnPUSpUu571UOE86o7O5hOVkFQBPwheN63GdoGSnp/2Ir8Hp3ptN4D0Z5o
ZPLp77B7S9H46VUIJAPTZ58HWzy9zA4GSTfFDwNm4T8uWPNw0ROECKFWm40vazk+bofN8c91mH5b
NIrPPzVDQM5XG04lXtPDntxhvX5mfy1pFzl9/Ko+TD6rBqO2dGtcCFppgk1m1Wb3gDlgWVUKvN7C
7Wvf87xmgm2wcg0cKPyqE4KVVYu+F0qd03nIR5Qj3Zp15wm1B7J5U4nsYAQUAlBuMj2xSqEJO04L
SFltu3j+NkllGxejY2HVEHnMcWhEx1oWswqes53xR+NqxNrS/pZOrEAPCzdbilFyadgDtfOQEo/O
oJEkERIoJRRn6cXSSacLIdmpQJ59sGIpuXo0kuURaRO8d3fOWsQjO0Gcl9EnaCF7hdMf0LigWbC8
EjmzCIVDa65pLPmv5OCw4/lp88egUZgACY+oyWGbkZooUQ2vNTC0C1GeLIrO9yjg3dk81unvTqqq
rZLNv2ys+s/gxK66OTFlSa4/+gshmOMF4kYCIMMXklar/MeaViewFb2YVsLT8QiJ5yHFnuAZ/CPb
pbC/HyOiaVMs97o8FFJ5/R8iN/tp01NUAgVucLu+tgOqOYdt3UnFM7r9nGBsU3z9mr3fD9dwcoDG
cZ3DvB3teZA2qWZzGF/rk3fZoH5lpNf2ufzJduYfpdUsHLbUqxiWTBQSsHKsnELtUakoo3Sd9+6e
usl8szynntYJ57HxG9gOMxalGIlUZqDEjfafob42X9KVoAFf0V9tyDiaoGjJLhqM0P+DZsSBfJQY
Cl7p/DDkI9hNztkE59zgNXTq8nM2wf5boUOVUzH/wqbQPcVf1IRqke/6L230lODDVVPVLpnankMK
1Hc+G6tiWgUqoAmyKJXm+dUmBj+/YC4Y+yj/mDjpHGOdlIPYyi9Fb6Tf9nCVYBSkjpETLPmxAfrT
kcmZgzvjgpGilhzW6Vv3JTyZhgbFwUckF1qCdnspPiw739u6gZW+wUWI9qve1Qi/60KWh92n2wyA
Po53vhWjyf2CVoknzQ77oUf3PVrPWaoFdpm8JdUQwM7Z9bPvhB8V0nnPPfDcnOnx5ZoPt/wcBj9s
GgmFIszl2Mr4wObnKn8AVUmVyV0P85euAAAtVrecYpXMHajkOKPsdAIlVEMV2DFSCPnQd5mMq7eL
7X3QS26c3wQZWNBtkK7WWZpE4k1EPTG6nnvClfVMmJUZ4fGhoJuAd25Mt2arEIi0ccdo9xJPjaBY
LSYvxDDBp7aXJNT/w6PPMRpUPnWvytIa9wXlr2aqtzCiEReHo0j+PCFdSNCqGHuQqpw51A85fBpn
pzIYKyw+XI/IoRoCNommuPs7Cav65uJ872YLMD2BMiY3T6TpTlbWh6HainjbQMiaKg/H0Dz+H37q
hYNldZ0pw+XgZ/Y0f39WBKPFYT3P8bqSyNAaEWhtd0KtokVHdymTv9ZAJaemyZgg34+fv0S/WqLQ
yiYUFvGfTONOcVLhj2QhwFQkFzjbn2s2P2QIuigKT1wYClu/l+IlMXSLoyO6EyWLlN1fk5hmCQtz
/AC37eZHYd63biGqKFMFdmcmOnuc6dd/hKIyEQF05ZxOIVF2h/HkI8sCoA7X7lGX8mqfyvnmQlzF
DaQ0KZwkkvjH0lJeNUUEofk1OEOwE5wfujUTezmbVvjZjQnqi/v1qUBLdps+MB0edRhSv/HhtnTe
/ApYpUl84JHLy+DvBDA1We6E/1fSfBSCZqyMGs/wUrvopOX4lbTfUNtIDYajOYdJjykRoVXhKnfW
+PCRyn9nHdvvf1gW4YK2R0zH4bR3JirNKFm4TqHVY/7Ch8Shq2PPTg1/+pBhXUlK1BuIsoNXFUev
DcoiB88MtUreblUXSwAXB7kWlkF5FGtkFOyPt93DL/AHjmkw3tPq0UWTljWNS6Rqm1N7ky9qQgBd
Y1ntX91DkJI+H+T33GbteeIQKgBsUGpY/ufsOXViIthVtP+wwXAZtF9bj111IRY4gBHX8E2vpsBw
eK9Oz/v/Vu7eoWNOFvaYnRSEdXbsnWGvPkVQBySqtwAJE1wQIe5Y3KXI2EZPJnE2X6ywwA11pYWQ
q1Udbbuco0XAEEkoiw+0CJEv7pIKeWMsZzy07WpyjgdwzSaMIpJQX4UkENMsm8viMdGywu1rWuKW
xxz32POD8GVQ6nofgcXlbL7grXDTbjlFvDrSby4wK+64oJ7KO+s5uId8DHUm8s3ecGjkNR2TGkJS
PyH8R3qRM8LLrMMG3D6vGDK47diw3xpxsY/WAuPWcS67RJ6PzgvWNj4Y0EkSI7rrrzdO58erphY2
MKOo1fdnkgIgMyReW+9Aoky6yJMp1y65vWQ2S5CvkhHLMS/YSG83OX0dCW91QMlW1bUU/Tg2naQp
/DqvcMOIUVYcGWysjWiRXLaxZozVlPBsRP0VhG+g6jz6OLhUMqxyEffxG/xz4kBJR5+mvjWN1X1W
91BblqvYwsbVAh7j9lXUDvhyO+dXWr47txfyYqJK628AYdi+1C04fVLsic/4b1xCnKy5qXhQQHCw
GOUgs1ZWFa4tH7Nsi5GxBx8JpdZ4unaahyyrXOXy5FucT++UzB6EoPt4snB7pHLFzrl2mEFn94vb
gQvehUmRbTz/LauscMjZ6CIvWqVWQoa1ogZDVFX6CMsB3yPzqRcinTe5zYmBwRe9bING0OYPP1mj
hXaFkvDjDXLl7il5FtBBaAfEXJb5FkAc+jBSXIOdaPi9jdwWt0brLg9n3pEgix/0wPZ/fuwt7wd7
V9SzhMSXJLNLuQAxK7H3MLcM6I9QblD6SqB7nl22czkQPUTp3M+AguAn1cy+VZ6WlmsZMIgNico7
5MxrAS2ChYHCT5Zbh/snIKi6u4NVm2DVEdVs9q+LIKworGe/NKzSNmmeRUMoTevHj+fL2spJu50b
Wyq9axQUi9uEjgrh6uek513Lr0L81T4yXCj3YsRSQUDOGopKZQAnp3UpHrz8FRkdja/Qda3L0g0X
0+iF8Sd9+jG2pJS2ldmRG/drIRnqoYxiVSyPGhvOw6m1WXHtT71eZHJNoeyOZHu8A46gc5KRntwO
DhamE1eeDoRrVky8l9A1Y10CuKpLsM4+QpQzmHDG4AddWZJCDRYSD9hcaBcI/rQ4C44arZR0paSk
VTM1378x0pytHfutdP+5rtcwVnpIBlVcCGc/TeNkrusZV+fbRGg16bfTTyZa791vQejpcqckSXvG
eKWa3OAcAecE4v82PZdhrER75He5Wno2GnaGIU5ho1K4eWfgqPeHzHOFDCeKMbWfkx8Rjh1RRheP
x5MvXqpxPAGXUZr4bwJrFCOqFz1WaNm5FPxqmlq3b/2Cnu4grAiWT3tX33OKlsIbQ4Pq4kUomx+s
vcdry6EGXU5dLpB+yfDw5OeYHEb0GA8lnXIcea6FkBq018kYfsMo9iTNmxYe8WI5rG6hEjkPrsTh
eMt+r2YNn1kaoVpmSLBRuk3hunI95KgTg8PUj94ndhdXn76hgcD1wPk7zBDbam3L5W9mG/Jpf7yO
t0qpDrPkeEsydJL4n2TjEk9ffC+1av3zoSXFqWeCFwzJl4oKLt2VJyBGXMw6j5iHP+wMSjyApRZb
dHxjhVW1PWErWYB6/o7XjYlot0Vd/vmWWNFm0QeCR9VsAQWNuzvooPXIgHs+0tzjLcH51Ghuq8Bt
yz5ArE+PGt5L1Uh9sAgFyc+xYFFHP6VhpFGtLSORymazaNlxmTqYDnmjLoKWZgUMiEtPkPsMkFrG
B+KoPCe/NAOn61aYL4o4rS1b9LG3cYjUYIx7sD34ajWlGChz77NX1MmKBdESmNa4t8iVKeEo/35t
YTadncqiHo5VVPUnVbzQmk1SU63GYiKz6pifbiKkvs/DwzFFKDXsOyPGDcRYSTjaZh6rqQh7UasV
O9B0Cs9Sgog5ieZ2Sif3j4kLMMG9f2OtbHbqGPM25V9DuID9fcHaUK20bjnJWbpRKeYemhKCTknX
lBlYDOnHqwsxxu9IcL5be02o6McsH5XGxZii1BVfJ7hqYBUspr7+zebocJGunxBsOQdoIDiqvSV9
3S/b2OvO3IIEXcB3kC0WEiLCicxKsrLfPiv8lJupED9fF8+tL+WMjluLjPWWOWHvbpC69i8NMp+1
LnZTzo2h94dVnasuSfZXMJ9d1jbaVEPQTK9R0e2DrK19qLg7RqwsPjv93qq0MNCE3BAVccyud/Eu
nm6uqYJEFMnIPCgT42oCZ6Q3yKcrQMlIoGgvmGWalEOVwQeqehF9x47TqZ+x9TQ+xnowPj+9j5/f
utWJlYis2wzvdYLpwMg4k8lyMWengUE7WrasX8DUfkqyVxeKeQhm/QwLq8S5n9uSlUFlnBKq4c2r
fgzu7FUPv+84jQznit/wyeuOBJxEaJxEGGXAcVbxM+ZGOnjfQAe4S+BskalJP/CeV8l9YRGflPU5
l7XvN6AcIdNlviXT4uEEgi2bbSeOYS9WFXQnX4CM9zi1ZAaoz1N20W8CcTqnh7TMtLFxXgUPu9kw
IFYkJlNSofWEGmMX3SGcRB8K4751Obp4ZndfOkQpKqBdWcjbzWnbrNn8l5NbvEkZeSnlaEbslFs+
HyfvDH6rjYS/0vUEoLU/0FVICNdLENc5bSCftuNp4L7WqX5uoLiChGS3msm0r++XVkDOkPJDmDsI
TLxvN8y7quZXkh8l3IbzKC2ODAfCW4ZeC51+pqGB8MJSgBQVIa+wr0awKdbBTZmux2bwAriY/YN8
rdBryrHNYHXwDKdcwH3JtqwF/GjJnHFcz6jNo79wO6fp6ceuvRT+9ySB9g666uAwfcwkpukBgeVZ
MNR1bHcLmUe4zmQMwVMrI9C8ChCITS6sYGxj55jpFQKKpLboFPACfU09FvOQchSK7Ckll7GdKGu4
0E8W9Qe2poAZnHpzMlh4tZzUritBXvmSI9w+509ESDwkcLM/XMrxAdbvCCpc+nIlwXGeDnC+tchT
JTJBYL1ltNsy12Vj705E2bADGhLnjpZrkmTyOS+fujqlwoSg/dctTZK9Gkqb1Zk8YnrpNept4Jzz
VQTX1x3fni5VcoX2bukiSe+sa2CJuDZUkpuCcM7/QWMsMEc8mAjk+gEQgHhz0QldLW935L5vGnY/
tkVFt/2L4Km/KIPXVANLOsMz/VxKBar5Ki9vX5hjrA5NvhzQ3xXTJW8AgTI0XTYlOCKZQyqM7l7+
xXUiIXu/+7sJOsVPqAs8Zoq4bJuJpYj8SmlzJUMUC3LSu5kb6zsP2X3puuIqmtAuVWZ/3+7Y7lGp
DRBPhlg9tY3NeY8EPrtuG9bwZIshnsF9CfsGxXQCiouaGaEoPGgSX6GF4RZfIi0a7wwj7T/h0zu7
iRoWfSUBVzMfwM+1OP8Mks3EExn5ahTvwstKSUrAmsEEP2Is7UcUQ0PD2Yq10ZumJKbwj6TYHrNZ
q3Nu88fJt0Cp2uRGyruR1LAm18MsQH74lEFFz2p1OGKCuIuv5N3quc8t0lrbVQMZ3Tb6JFzyr5MV
21iBrHze1jZYq0Z/WA7sVVbPQT1JHDYsqvepwmUVogdHP9S+/rTbYR84v5UObdvqgWDYsDYGTBiU
nQ/yQJicDoHWRSHwMlQhHaakYygScVD7NCTSz4fsaeTPEA1yTqnZyAlfxTMVtv39uBNfX4aRIW/6
cS1Cy3fJn78sEg6/nDfgTQjUtLJM4NcbDAoKSt13+PVr1YU/J63fyG1Ki5PIH3bgtBIvZUCfAn7T
mxZKIrEVmyp8yvUSgGoi/bQemjm28ebnZTdrdlzEATpyPCEwM0YhjX25ssuqbr93RC8y8PrU+mUD
zLLkoRziE6YMRtdqKWYC8XZf44YidGycOjPyjZIfB7mrpFHUsce6gucsCZ0gFVp3jvzYuZoPjFys
0A8uZ+tD+rF25lPt95vFNEr39fYF/vJOFA9GFE0rBzmN6IhIU6hoGMnxBGxb/QApesPSWVcX/339
BM1px1aCaoTSOiuVuex89cblfKHLnksFUHTKHFaSvOl+v/jyt0drRhhuOpphV91WdpMbAfG1NAiQ
/K9KW8Ooj8bQernACHZtfYF+Z5eS/0fYiDQM/C0jR13O3/KXNQ1Lr/2rOJFW6c7RUfteyUt2g46g
lK0cmipTBHLfg2jKXgKwXlrSQ54Z0CfKbaowqunnBPF8VP0GaYnU+/Fk1CAjKOqsXdozDjdqeAGk
meVCCS8i+BvQYB2T1Cg6/sOvd3p72sGNwONSWWW9GGpYBDdoU5+PAkftfJ+pWbr+HiOqsTce9riA
Da9hC7o+JgY2eFnolyVNvk9Cwk44c6Fz7n67D91An5mMZ4gzmNxVukkHR/q03k6pVbX/hzqxc4dq
kFmNcRzT0/O4Sjyk4YIyxK1csKZccLG0af2oE9/AKtEUvhTX+dRRApX7xevm6vNy9amTTOBvAJRv
9dXPkkNLt1Oiz2KeetAjGRLCnfYvqPLRz/vx85oLC+HWMGoGwf0a5hSJtaQ3SSoR4QHTzei1wHI1
ac/x904+ZvB1hG3Q+TlmfyLsi7Fl9xRND0FDA0y2KT4BCPVkUXqrv2yuTCfvFqv6WMujmbRD+tsR
Xc4FPf5FJ8xF+6+IhYm3RsHw9+WEqrliLaE9lCPXwyKkSWoAZJspcNoWU51xFeTFaTxT82Th3br2
dOczfMcYN5UQwNybsiDCwSprOWvVEZEcVBCESS8e30GENFFylWoGuqpZ14zGso/9A/uBtJfXKeOu
vSFdYI4Vmu4wslbezLKPCCDbSnbtui5/LwMWQu+C9UHEGBsXUQ1XQiFrdpx9dfEm5McvxSTyrtn4
Kw8sUYYnQbBhVfLSQleKH0z0qzMUrc21IbP4r2T0q0zy8gjN2inezU0BHd6iMfmVHNOl4RtjSw0D
p7ZBQqc/YRgOHQ5MWHeppG+VJUymMUD9Wwfy9vCxiIIA6J1PuaYOLBlTO8/SlZ5SnOxMVuJbHGtH
heVcQ0IBUFV3yJMlrrQ7Nzh74Pf0x1uMukeFzo/xS2P/Vv32f3B17drZlt37tK+QLNy2Wk1zoUYy
j52Mbp0G9TpjWvsAAL8ImH+8ZciJex6TyaOriggVZeXEvvsoTodLz/tEVFfURtB3E2j6TgjaviR1
nbFFslcLETC97mw1oJjgYgLWwFdQdJjsBY/CoFIS27Ll+OSVbSG/HWrEs7sedq540NMXeVzijmJC
15HQPtznh8sA3MACggy8MWw8whptf9SY87f43zWpTheSfZideEoaQ7iEiVRdBcspO8kntkFV0CHv
jBNSHT63jVrwi4+ogGNzSnc/7+BZz+eLGSPzH4VVYllhu7qx82Uxo5oKIbHTqFnQUXAIcYEYuq+t
mSEvCtmLzWjEoAqkMT0PsfKQH0IqAdEV01BywYJzC3gfGshwZ+OGSDYbwvmtxJKjxaS/cA2DRhsE
ai3Fq4iyCUYXiljsb0uwfe6Rj3AfsV8mZxRhwu9Y6kkkNYq3eyHdSVTJlewBhamgZ05kVaYnBwyq
ksdFKFTc2WJIYCLixlWli/kSCnhdjsRy7nN1DWwmFVp7fR3RbJMFbjmGulM7u4nYadFlNkFPOjnO
x74BBnUr7oHbHy6q9XrcwH4KEEIrG+2j+4dTLoHPI9ER66EZcTG6MnqMgD2TGMmcXF7kFGVAumqp
tkcJUAKDqAu58gI4XkgeOchRsKD4dl+S4um7u/sVhaebCOAlqHrCwk0I95I6u/yiOAvxqzYcbnMv
2JHPEIcd241lILtsLKwiKr5y6OG67Z3FYXUo2rc3Et3ZkF5oHcGSKJ8juWumagjCUdjfPptxpv1x
A+zxVAoInxGaDSnit0whQwBGh58c6NCFI1ZFAmH3nHF7JbfqNspCZu0GkgSDXzxcrGD6D3xpz0Kx
FdfVJjYtJI2MAjuyJBM/eYuDVBB/qGRasOXIRN3a1nX+e1RVKqDO7/mxP9y+NTzF/DYX+ozPfNvp
/n6nrPa2LVZaHWVokxV1mkl90I2aaaQKYoLUsF6zVMyA7kL/XLP9isXKOuZF7uNq7w8aa7yXbN6n
Y1XI9RCTYx2qQt1Y6p3G1iQMl35DzQiMfjuGw/1j5aXOdTlVuobYNT7dAA3wjqtqwpHBciobv8lP
DnqGKHs55vCOzrvpkS/7RHVxZRVbfqp7F/10BPnGA9Y7ASuSH4naJ1R454jKyByWwEwKbWjd30YI
J2OVg4tkEWeS8/hphcXLKVtoBKjvYE0AoLOrhY1rb2cmVnTH7dNZaiq0Yq3OI4AeZG/zP5sXHmgw
yhizRJOqszj3YxpKsToyrnVv81rucYIlUo7D+gK4Y/Gg753WZ+sBvdt1YT19cYQCJooJ0ieBykNF
ogdmWwFQClOnGdZHsps1kf+8pklP3imMEGP2aGLIXL9In4OVuf+32RlCKu4CfXIPiQJv7HNNV5z7
c9lnxBH99UUaty9GPhaBHOLFp8kAqYL46JWd/lqhI9y0DfrYu7Di0VnPWHZWSmEekfUKXfH5QZAE
s84Q5gp/++NzhIFSs+Sen+Kqj6MKGs5JcLzqFEuKYB4FozmltXEDqUCd+q28Mmz2/0efQrYv27NG
3tKICQf6dMiJ7XogFMdF+EMnglDXgCWvFbKeQnkZeaGQIqL6xc1vSkCkkDRv69PfIScYVJXfXsoC
ppbgJg41fLU+skd6L3jhl+Z1ZpXBuH5wE1ej1nAH+1goA38o8yw//CyCP2gSyb9Rx3RS4jB8la9O
2kv5Zt7BuB5xEDRx1irbrWXtaGhpU/QV0gxNpwmdHsjSK5Q0Dv9xOrEoUvIiJEuacqIpbD+Er5Oc
gBNgr3uRjf0yYDP7EfkWzhhTTknof3d2HQ0jZRjX66WDAy6D1gt+PwF/fVB9ixbb2d5UIVkhWmvb
8/DXwPxHMVUyT0sIDV+migxk25Nij0pJGbE4NIYhezmFHC53dKmA7rJqXZeO9+ZohKtGunI2cvcZ
nvAiHVlivo0gBIetihJgY47YBm/E82oSqio05Y7cUJ5k7hP/e3182THYSiOn1Ki+0AfztNYf6EbJ
rY8nHBWwi5uOdRnfp1DqRb9VYp4JwUPOYpp7PXLXdE17Awg1SoRTIu2lMYjdIkxQocTJMnYYNNmc
/bGv4TwLd6SfemVn954/B+gSqTZ3asM/5grNhVoigfSSCLqCzYzTBYt8nfNhfoYtUdhgpaBIF/QA
8d22pKk9kcejEM50E17QqkiR5p9iTjliH7m7AHdrToA7WDECAy0asWVT0rQzP5DgglngGMWQLcC6
tlvzq9X5JJcDDQeFih+BRXgQcbrX0wSJKFp+PQVrWix1K//3ImqBCtN5VQbQU2jy+61NuIrQrsaE
o5VP0cq1vkHlSypr5ZZFEmYQtqVaEowWueYWFm2k3zgWFWU4EWvprTSDB4ANW2LkrWGJWV7cR7OF
CN0l8rqh8WoljQgmjCXDGbtcmAzNABe7aqfwOF+KIWu5Uefil890NHt4WzkgdD1HDsSZv9aO11C/
oEXQPm/eVmjm2UJoH/n/AvEBplpiVWD8A9hVHYS1Pe9zOyPm4pwn85ovCawBfNOmRaW/tix/fqUQ
zlCQCWZ2IFh3ctrxK3vu8aYfz7i5/7+hlJmDZ8CDXZ5H4sRf0qIO/asEKqSggnQW9HDk/1VKF9/s
kLJLoTRCLLP6djqVbY17xJOJxW3Vc9IMok1kjP8tw2+uX6kfwzN3WmLcvAt3sqvsL9ai0J3d8Ra7
h3wjsaEzqJCrkkUh03mwzMJgrKa/zj+LKAaIj/NwDNz/1sBrPboyKc+LLNWUJzRns3iTnzVIWyKy
hNRJFGET1+vz9KtSw5ByyV6OUSlKLF0YXn3gv9t1b0wqDt19Xuti9Ydkdzn7zWMWkGLFGUWSRPNY
D/jCOm4IZq+QC3gyiEofLsMjELCpTPnFolejrHpDmscyXsFkfqnySLkjofCsKASLUe3ABO7AHqQ7
sslj/EasIrgNXboItuZqPvlzU6ujk6RSvGOnIkDiWJny190diBmUU9Xp0l0lnKpEiTkvIzuQulPB
hyh998trGZKL2ZZFmtSdOE/n7lcatSvISHcsNagf/emGKempB1UEtop1R0yX+pYXgWQ6aldD79gU
FQV3k14X3Psw0OxYvP17ho4XnxhcOdNxspMGrJeEEN6ENCksZXfhZTe1jlDQaNHAlOaLLIxFJcxE
0EBhGX22QtXWwNIYj6MRK9lYHon3T0qpa6ZdYox44pRszx/6vTJkJakK4i8vnffLYu5phM3WzkfU
l5mf2kK3cJEoWWkxScCsAlFK4uquiLVqTX0NatcN7mROfM4jRS9krNMv4ijaIsqF2WDyTytUWXTo
qNESx9dbcZmbxzK6mFdgcfGRW3eCTa+ui/QkKYnRKCXBDXeykSkmKE6JQbhlH/AsrZ8zi2kT5X1H
f038EOf3weBqZX04Oa8vGutrlOgulnh+LbNsOvGgh1LALnYaK+VYxKr07cTpMkJC1fzadFrB7c/N
11aaGC1Psy6A1H2tYLlcSPtNQjUeJ72GAIiTfgsUCJQxGD5lkFF+TPneHrfHLUhhh+gkCoM7FPnE
1MKoxONd1ynXdREIJsyYLO5JrNoJScWuu5I70tWKKklfFeMy0VsPyyZV+aCPb2VIiU+JxoyF5ICR
31GuEGIRAE2PYGinmxGazziNmmh4T1+sqBjsESnEXJ8GV4metFDO8kzgW/BjhJJKGJ9E4b4eRRoa
TINHVPZYbhgYU4q4+Dp/8Uo/mpwaMqIKDMq6f3Z2hgXwiFAjF9h+PjTWPYFa1wK9AKX5tL1AoLJ4
vvZCzahGpaw4KuE2yKwbQb76jdiPJWgxRWLD7GSnoUGV2GGL2cy5CBkGG+/fJhpvXUp/aiK66LfD
XR7zJujE7tD4nqsO9Oei6iW1RlRS3aHM7OhnhVDrnh2Aaq5iSuTemZOrA4cvNQTOw7MEBxLILexb
5QR1yI38s0LP71kyzqliXXLZsnEKfTrzp22DblB3sZfzz5pMhmlT7beToHhJdixsRWucUv4ZpRHq
W2iwgGE5Kyigbl3AwKalsfgt8bpAz59roHiwsIeq7S1FL1iubPVG4Z2MalDYhm2dCtilyCfSe7B3
j6vD5QwpCX5/XQLzIok97YytqvEJqWPnrylpRCcKC+DzYKTXT7ohOfyXE/Q3P/aCi0UOfFfowrhi
mObaRQxg08aoB69L81zaIVlyEiqiXVoYeYUWq10fvWelbu5OITEUEuuWXfpjuHR5vY9w0aDbnm+G
i69Y8gh6L1nhi2dIWzhO0TsPT1GarGry6D4UupCwWZkl5elEJWB3v4CsWPtIuAOfOb/UQo4tCWe2
C26EfckfKaitlUUcz+NXAr53MSPg8TGhdzpXoTkkeqUWskwmLlKHfHYJXoAMCNi0h8GRb74AZWYx
aswiGieFIMl7nGd+XFysYSf9AqmZZ+r+bVEnz0vkkBVhzMGuHNy9A6DcawUpoVWE4iypyTqHmY0t
BWXv/4dUUwVTZebZ6g/Y2mwT0i52UCYSUMhJho0n7XunUOE5V/6715IsNsfF9ByMUJEHxBYU2rTs
j+WvON/z/Lf/3SbKn/skjdlEydAaFKyZl6qD+AEgK70Dt1VENp35AWydlZ/Qar1nPRnjOnrzQiYR
cSpHSvBvxWxzgE5tPLgzfieaLexQMv5zaGRfXLfHFiTfD4FDyUkMpVH6rWA6KndHcuwPbsbYsicg
U539TDrTIMwSzKlAaT58fZEaVX56cH4Utgfe9mzKFlvVqJu9oZHPmqP7CqpN0xtCwaq89Dv8F23/
tnvyho9imJBZosEumqbD4pCpXONf+BbqWxtSpblnsx0hIDaOGhb4Oeqd7TxCVe1B2vjVgcueBlYS
09idO6fG8731m6rKIEI01iSmWAN8vj2lnxr0fExltyupmQNlRZiFSIGNVAxknGY9LT8HHX/SdMCR
IHVO4P4jpKITF+A/6ex/p9+pnDYRlbzl0EH84Y4wodHhLdJJHYegwIwFl8hb+0EGPljx23iaOfwA
nhuaoM3+e67uH+rr4+hsjPWJzMPIQKuUU5pY2/z60LL863GB+7151jyVgE6N1wicR3J4td8kQ32m
eGFILBCqJmCU6WqqpoFTiNBTq1BnmHrTOT3CCp2CdXIHsnIU/iV23yjBeCSF8FN5tG/LzbrDjXt5
N51eSsG3m1lla8o874ctsnoZ5uwf0L8Exb/F62Cq6mksSeKTItjwpLIj/r7d1vQqvyi/zfx8N1WQ
54JjWetRFAQVwhFny9JQ2pevNR3rAAYc3FOkQSFuHKMV9+c8Z4e92qwjA9a9vBe7U2sYEgTfjrlB
UBm3GUFkEFFMOnlr2skYUS5lvp8Yseul1S97R4PS+gPsWGXX0p3UlorS2R76Ya21f3Hx7eNj4hFd
ah2PicHIleN9xfgHXDHERKCo6ENIwrxelwroa3rzQHaSSipd+boHz56N/KpBd8AW9Bl3F2bvo/gA
nPtOA9ZPqYP7XK8r85n1VYYJFpRUHr/gxLF35GC6+iwD2KaDo+xof1/Id6H9L2xg/tYFVKPigHjS
+Xle3D9Ah68Gchkts6EY2qsBKRCNLYGZEac1cIA0C3JkCPF/zX3zDs1JRqKJQcOil+j4+95Lgrxe
nwRaygmD98BQhDzrJ/qEbt8l7FEOMMwKtVAvI7XoXnrUBnDW2aoSxg69ip7Xf0nYYD9XY8PJhczj
AHmMJMrJ9mjNNH5ZZyK946kMzA3zaE+Wq2nXhGWRAqyHvJXH72ogdwnaCkpVvcoLCGgoyczGreaC
4yHWjq72f49GJNzuTqFvhcr3k0yNVvdOc3pmcqXyo0Bx/REUPBNk0TOHLHyrUFGpyMLMGADShMzy
tundGIJ5LvtLV01JQYaZ9ishkAi/C57QUS6PPHCnM2n8KompFfhx4fInO7SBPmPxLzemt7rklUa1
L3zE8FdDjxN/yowCiOtWVhqmC0GXEBtOvl4C8ghPPOgJYRllolo6RXdbuXPZI/t3KreSsDxJOoUW
1BMhn8LtQ1cAC7WKiffckJMS3i0uBr2VSECKZy5BngkH5BQwCaFxiQp9tg97QaMv09iPb5XXFvc6
nyfxiAnhrDrVfPMjnFjxYvPdM5h/YpKUFNPe1HXL3EeLFpi2q7BhJTnlHKiz1y3XYqUGOcbVHCNt
sqVB8vIpPaUwxFhaU6Z3gwIjNW5h+ys5Q6OBZaYg2fu0w2Bp3r5g2sokJTPRRS9L6fYeazpR98i1
HtSzzkwUNUjE7Gq5TjL2WZq7wLuL/9yeOmYECWmLfAV9V0KbQe8BOrCtXKIBtLFr5KT7RpNz+7m4
Kjg/DwIImKExpe3aHnA7z7zrOeQgnt58zXV7ySudW8mCeIRP+6iv8qL93XRGkRvmNYztn5pttkJ/
hG1RqyQ8Dd7L4TcE0PDGdPTJXMbgwX2KOTIm6/l4RrtzhhT0EyWX0UVnQ17HrOp31pdbsQEDYbMM
OnvcRSUJo/WTJ19gBMbgrhL6/G/5BN5AdYQdjf30v3tYojlm7sHbwzp+qEFheJ4DSU8La3xPhBur
thW5EM1tMTRqNsQUPf4lkEXevcCx7g28qMmG0RkzmO78l4sw3rcuwNxO9dP5NByeozNYUulcuPzp
7S1ho/on59sVKSJz3W1YQZ6GneU3vZYyPQp2lHryGcBpgx00pF8gc1D1ZN4ujOPX+cYpXxEhxVa6
rQQCDXj0WEVJ+NmdQlUWvRD78DKWDbONv4F6Axx/34xdk6y6j+bbs0r9KCcSA/S3sz+SRmKLjMRB
v+Y95ovX3xbB3cKRPuxMtuhSDc7mV2umsJt2IYfw4NSA8+5vRWWGgLCh+v0dqrC9CuZ0/YxNjdbn
kDac2+FEAb+I2FvM5K947r9aAFHjlMjhX3EhbBgEg5fxcdXCcXC28XrLWq/HqoB+5oOGXHw0yQar
TBpHU46BUoQdH+hGoZcgGvbG4N39fyTvaDFVp5edYCydF71+v47M7dj9OHaOMOEcs9s/Lbt3ahsM
q59ce10Spt1IdGiyJ9wPd4fdeqxgaPCgJPZ1e8JIpFyHrjcmoRn3YUqxh+Qt+y5v4CyEojS8UCqi
AkUxA0ZFhAQDFQXJSQ2zAujsaWJjZ5PIQaDTNTjGNoF2dRVTWpId++sbyDkdgr8rzybsuuIPf2BM
DVE1GD1WskcSAFqQefHacGLavPN3/ut0KrckOjoW20fICMtApsWeikltoO3LSnp8/t2z5AJO4WcW
SsiyM9Lbd5gjeyiv6ibyOuqorPc0B4QKkicL9TbSt2bBWKpUmMkyzmQ0x+K1/R51VU4H1hLopI6V
mDP6mdvA2IvNNtgYEqpFQ2nzgrYla7b50pJFZdeGhQmKal504mIel56kD8EgPXWqyI+YJFhzphrN
strT6m7lrzvLUm3Bfwv76MecTXO6nEBrbpDYLWsi2SMy8leWGFZTJZg0vwQrkkQzwuolkw1VJ3bK
j8FrPL7bh/4qIFH8bgQI8bXt4GNvdLkJb8jOc49WrS6JWfF5BPBmXwuZyeZ7SFGx2uf3Ep5coRHy
39AZQWeIB0bLjJZyPPmYqnN27nzEa22AwSpMntU3n5TU4XzvHm0de4ZFMkufxkAaAj4zAXdoLUJM
yj7+5cPIh3DWduvnOMckwED41Kd1JS0B0dHvd0g+oCktBit0Ln542wW+KPGMXBTJ6IUniAlybkYU
73qv7iXmiIKS7zjnwAFv6G6nsOxmT45C8cd4cGOULX7M/ON2nEd6FGh4MXDsxhdU0NpQ7e7fxaUY
KgkYOkCgy1WOb690XIRw0QcBdMnf0hvXZABi/AbO3FeCPKxfS7zKFPByJugqF6SXLExjKpiLVqcy
6nGIIlwS1Q7Asj5w0nDsfbe+zQzywKbkfIpuyggQxb4rMNfUOA/RnvS87xcW3UAwmAUnrwQIvWHM
OxPK7ZEIUaHh6VCT/BcTAgIgcwrFxmF5uUkECd9OqHtBewIExeRy19XOsyU1Qa3thgnU0e0tnnC9
D4ByVSvuMTZLc4Yd5Gb36WYxysmYiKumHbnTgwj6Jedf+UUoCp2T9IbptGs+9bW1Xjg7gTQER1Yp
JKHxoHOuA9WcapQ7oVWtt4xvj2K4j4ay9WsOI0JJOgGfWGTGplP8lWD2cxY8uyl2wG/yR51HZxuD
nt4hxPNlxsI9585+BmACGr6bOy96zi5EbilTLE0nFKLusJTUrjVRVcAOtJtLYggTkUSUFGIa6X/Q
//AbchKhqild7ItNI0pKkZvUyryqNmeuCvL/TU6wCda448Q15e42fjts45GEhGn0710NLsFKzWQ4
85X2Dua/8Fwh+CHKoi20ZG9fZGK2sujzvdSwOzU5jk7M8+sEhTPQv8xjkcVRhu5XJQ3V9+WR5Mm0
l5FxHxZDUdayIVudnt+kON4FkxnXEpfCMjorqRrJ20+1rEpAJBI75BlhBqNE82VmnVfRNs+h+1V9
B/oUZbXG/gGK+nry3Q+ZHWfstPFrrSh2b2t811z4ATS8Py1e+54TKwCrqkljgGSlicmaUB58kVjb
ytatnFTq1oZV9EPSCeHCaqbMU27Kn8iNWnK9Slnr4Y8BloGd47XoqUYystvYqlRPHDICDmRCjxmW
qYFImZoyx+zpWdUgFRwSp964PmXiy6rUz5poIkJ5LDdXbR6Zp46qp4UKLSjoT2nVaJDBbrdU5Wfo
PYHEhiGBl84XGnwt1J2TKwsV20iyptEnPejLPQjWOcMtlmK5YWo85aBDFaneN/fhx6Xfaq2ud5JY
hmR6l8dNyw2bD42a1or3t5oMZdHzuyYQL8+Vp4TtdmEvIBM0YzhAceTvtgjmOG5eK8pSPmtL/TDM
V1Bm7jrL49/RnbpOjti8qI3prQxfL7BmMbj6v83MLW2A+hA1IfbrrJalYPig6khar6BwThlNW+NS
mIDzIufzzFSFpaXpyzSn3NzN1PEimsCLnTX8dRLkLyn7TtDPjVTOqD8J07S1mUyQKbEQbEe2jEFC
GhmFKLKW1slLixs2oyER8xVPRdNLx9n17Hl7iJpoTQGXqaVDAT+dS9MoqOY02nnaNVRT4eWcmwCb
P+sI8rQAqRcxLmu8HyuAlvWgJvBN0FUYjnTraIMgPUvE+oiPhFIosgv1y0NBbpNUTkk3cRhl3ihf
FcrDCDNA5wxeqOl278dxgTurDFO474uYjBAgBxRe5VqLwmR6U0sVbSQbVEkltxv0ggKdJiycOzvz
rVGEom2Y9awDFysMa827J7p51DdBKpwHNaWX5PMJJGHqMb2TQSTZQQI1ryfpNXblzpJCZAJNRRHp
zSTLP325lHh5Ii02mTIm1LdGeG3IzNAfgv42AlS0K5xHz38fla3mJ42k/BsHwjCoG4DVAUNmDk/S
YcTv48vsKzMS12w7950tDYSuiCZEo24ZakpSdU0tMiX93zvGTzQ7ZfTRcopau3JC6dfeQ9URqEOE
2kQ+YamxCyUGbwUPYf2QNqYpsx6ymxbhD9yv9sW14NN/STS56zuAJAGWWQB3TT6mprG9hOaym9bq
EC3yFmzClKcKiy7Gwj4vhUre4W1MPuA7Jao4xy9aRQ4QW/OJk0qxMWPZP2CC1PfMrIkm5nahRDeu
yFY5PkX+ZNDsqpRV7rvdSKNWoMgtudbyLAv4LNIHF0QUDpJYOa2pXeEXnEnt44pTtJa92s7DmtR0
1J08TilJZkpl+9Kt8NlkKzfLLPGhTciZMSkwNhbNjBMfwuOvO86f8ka+k68oSqghiVhNXl0drKF9
mkXEZ+8RYMeElv8OCrZ+qBqtA6alpF09WFwb4lS2tyt6FFtkspLY3SzdkiVIYIdvMQGmdFu2P+lS
v4dk+d5o/Va7l0O94Oss4JmpwpdUjnlaxPySF6OIUs2SRs9wfh/e4awSpSgyupjU7B11Qutfjt8q
8XdZn6NY00xV6QN3qjJlm8sw5n2LjQCVYucIw73y0sgUEcFFsrk1ifQGnLdEt8fFG4Q7KL0UQaLO
GJhDm6JEl3TADrmpQ2xTSRodpqPcvQEZadPnQ/F0YZORBrBX0jekcYtxqYcHPtevUIJKGux5I08o
URARVSdxedfppmew5z1KGf/yrmkZAwmHEs4FKN6m1Oo1LDIdYTVsnCvzqMxPp7SIvuRqlBGscPB1
DhIUTPGu0Wu7qeVZkKlOC4Ug0q6lzMzDr/gjjbzb6nl3S6Zl0JBYlDwU+MnU4GcufG1YfCNfj8TE
fAlh+zJIMtccvj/nxHXfn8RAT7n68/X6UT0o57FVWxevM7JYLcDlhH44wvxP9IZxmFxLBZefoYFf
PEU3oLb/WwLVXth5wulqbaf9B3cAughMjtrGHVtA0rTXshpZnN9TMqSj/IZIMtzDg7vYy9GTbUxj
3JkEHGqUtN6l4ha20CxH7I9U8ZGt8JQrgXNMx1+KLsqFOfY38mBLy1OwAo9zWr5mX1CCApPEunM+
K4Q01d5wRx/6+sD0rdfUx9FzJ8YbTSey3sMhEHJ723Bp1s2U9vHWxoyHPjF9pCKMw85J/l3SCKWH
81ygCWuHf+znyLry62bK9gmtlFwWuMclRTLspGJhAJmc6ck7h1e9WIRnaggZruugLTCRgQBZ8AQp
efqwhM6ARXXGjfbdpxyha3/evQ0ZX2aE6QgMruPOif9g9ajukUxZa3dl9oot85gJa2zf6ptoimj3
l2v1+sEERq5B7ySefii9+ESOoeZ7njvbPX/v1o0lsiRBJhSEUqEkj8g0Z1pSqNuAdqEEIfYA1S7i
ZnoSCzzZdOfE4AIE59bOM29tcjpwszFtW5/Vo0LF7fLaQaEaS57IOVcBPY8i8QZC5St1nSyZDA8I
LWnaFfJ4/un0cvmcJ4N+tLs8vA9P25951ZIIqUfOG9u+14w94uQQZ1lYLs+bv9BQSBuLWLtlC/he
qh5SxLtqaTyn3fQ6YPJ3RTl+gvxxidGt2aZrvDP0FctdPFecwMI8gA+Vj0fgfAPDxTi/SALwzfz4
7raGQueWU6q9jIGj1BnW3TQ9baTBRKDJVqawnNnlUPWDu8XHsdw7e1juNOkWeiRbyk3quYE/4Yv9
r1Bcj5rLiQmUecdDp7f63JTVLi1Xy4U++mK4OZ9eatmBs+dev5bCEAwGetaO7Jrncnbx9tMW8+39
bNALVQndJPxAeFMN9MhH+2Z3Yn8jRRdYzZKsKqTo4ZFNaYlEG4flJu4kjPCC6HxdLaCTduXhnmFW
ASM/HOzlL/l0BM1M9p2YEOQzs9bWbHVYLVhVmGGm0jluUjcCKBf+V5mhyHxInIWzn8TyspVd4OE3
YqyZ4p864G4Yvxa68jkgc3KfGlxgMrfayKPAqBL4b7q489RmeOJz/0sKRIKOBesuqA0/cIHIddV0
wAP2DFwHGaloFv/3rnnmGwKBZbyHCItdePnNP7IIh/m1ojo8K4ABG7e6faDVd+J/DMTq2OErfBSU
tebHTHn5yQvVAjLeUnhJ5+QYkBE6z429uZC5ARCblMv4RK2fFt3500qGW7nWzxyJybNeae3X0Wx+
C7DA1ThC8T9Pvz4/dVHbtCEQ81omV8Px5fSVsBL10dVWK0a9dJCTrEXDRvQNx/Jdk8nEQ3RkZ6xx
Js9kMA3KUR/nk18gW4ehkanvr4wA2ftH31zR/kl5wUdAUhwTHCnWHHFmOHGrQqxIrd7aMVRcZHv/
0wcHXcLdPIbBXtPAVpPmdn3RiSLvpkQDbrCYgkzvSxNQXDt1n3lh+bE1VCU4cYYsfBFGMzOsG4DG
48XqJ53rTJ0BNs/Qnq/Xy8oDIATeMu5S+CEcVfajdM8ydM1LKt1vdZLp3WZiJ/msDhQj0Ok3fBc8
5NVH9o8wPQnlJpM3Nzoo6TH/aBV5Z0IKMhNgxU9Mz2H8ibx1wdhMsHE7ni8pHmGwPHUroS3jN6E6
NXETh8TVAmcxt4SCC4xOdtdUtzf1CAtfzHUt1CSEyOFC2Dq04xffcrm7BOJL4lqWNfIQrml7L3r2
/KS4akaC01rLuwvENnG95VNSfK7b0odH4GFVNLHYXs06/C2oIRa4VaaHV8gjT+ByVWgegEwXhbCX
zfzqMjK6azkpLh7Ftsy5/VYwHvuhSNdC9ut0CfRkNqSkV1ELgeGcGT+23XM/RA8gy+LK96d7AiHp
v16DaA7/nr6VWoPqcYZmKQ4L40G7Foncnf04xwf9H4BtMSZcXzAhWIFzx3QZn5MXFX7mW0aJOZHX
hl0d/a63byURdUMg3Xr7HOdLmheKCG8Y4K19M9pmp3YkXnOKVChzF2K8zEfpS4BjSjpYnSQm9Dz4
4cDRqVK9QqZCkrj1ntmZtv8a4BErBnvrdN37NpgCYfMXG57HLDu3HAFJfVdyHPAdHAUiTf4zD5PT
9VL1fJAHjw9v1HZuAPovDfjSh4DRQ9Aq1nnNZMfm8R+xR8DnPte0jQO9hr7zxrjF0Pv5i873p5dp
/S5ZpFa99aK004NaoPum6kSnhchweTg2XdUsuelNDUzAQnc6nGfMO2JVFCCQuHWEf2+DJsBssluz
CtU+8KpBzGccq22w8I1zGWIR9LQwGpDfzwJ3oVmNjVB4wD+WXP/mmxPq3w8VlXOhRSHN4KQYh/do
LE676WRUVvpdS2ErtSsURJ44W8LOX48Jm9EGGVijx7ghwZP3AkDJ4gglCK8ru5BgfagfLUqzqjHv
O92+oVFgGvH1ee4/SkUZPDYfUjsmsBNH4NHQyPBbUPoWG2qV66bNjIsR4GOJAJHZrpWcZeOJ5/O+
DT8pRcpBQXfzcyWzKwacnFks2vDAB3hgLcvK+qmA3PEdrXlcg1yxhKuTrIafx94Ff5Y2+5a54iT1
y3n8TvkMGSLRu2NaVh3m5fbtyOtNCYoBAwBqUq0ConwAOTskqqQucneRcAxIOCrLnz+eLrOc0kO0
jVSItE34/cHFrH87avgdgqXSt12uGk7SQi1TKd+FcZ1R+kcaEOKAMtOzOm/+h3E5uabZHOYDlElp
h5+Me59TtZJq2Ys+Q2Bu43P7Kio93vMC4E7Z6qMtLlpT92WEIkROfZccrcbgAu4hVSFMGmYkIw08
2wtDKieJsctvw5tyDxn5j4l3p99BZQn5X/7Y1sYbnco2h7Mi34nrA5ARCvJ1wsDVsR+EJkacEohj
uqZXETpXWBkGu+3UDph7qzsIkQjl4I/XxTyuyaDvX6RTXO8NsTy5Yit9DY9lpTO1Trr6EOsBaVBj
2oWsCZsKrgEfcEn6xaQKMJkwO4WUqdVGHbHrlCq01uC7Pl/qyzwMi+D63X5ii3m6+SdcVyqzKO+h
x074jkKNaMI1RZRHYuXFvg6BJjqTcmCMW5jTfrD4XaWOQDOvW6+TUFiYn40z0fTRCDlXHnFPvXLV
T67wfDZ3lkw4L9OOFjoce+/bYbPgKxnzUMg5qCcJPF2kvtbiIyb0zplAlnZDt0IDMMqlEooOdb86
NHHnAl2zg8ag7q7EzfpRkQGqc7T/DuStezfokpPmQbhGfZZyY1pFNfEiyA8bYw5Q59bMxVfi3TIf
NhILYryihJxCA/EevIeNihoAB3DmsZ4GQRFvHxcXpRaQq8fUyhdtrHF7O+YX8FWaC+pVuB2Fe/Hs
9ANDTvtJN8puhCPo2xkck3vOJZ6CqUXqdBm5J6npsjSOiP3BOGCQA/KyVHGkxwwDAGH50Sz/BVzN
K0z5Zb9LihTONn7e1fw6ZG4IlidimI2IMZFqQcNY0CP6l0z78czG2k6qyvVdrtNi5ta4ZLA7qjfZ
1C4tcAh1YkpEdm911/pUhU/74c0y0iJBrWgV66wTK2KeqtFin+kJ/aSdKlzV+sVN2mqOMnIFny7B
kNqFRc+ztHIpXRYbL9+drVYXrOKwEZs96e2xViSai89XA+JrIK8tX3+q93lfEDIduaMJ6zv8/OE/
5LFFKtu89LwEFz3d2xmCkYFS9RovRduvIoKp4jg/IUKNiQaeDv/6+kzxGdM9sqmDFU+R8SiW093G
RaVbfMfNMBn2OPx/t/L35OoN4iyUbiglNACEWvyCpMzvBulfkcxqK26Vx5TTBq0n5m5eV/8EyAOE
r4IgNT7HZFehibdWrQQeUcVycbJF3dosjB8/0xHcsPBs8EwwZfiQtY/SNjIiDW1AVFfqeAbfMJzI
sVcQPaqq0ict3Fc2VC9GfU69JUAs02DPmBrl01QZG2QXm9gaNjrlRBmhZpoCVCgxEcp0q6Wu97OC
T4C8gnLPHKNWe3d/VcuYz15eGmx3XC4SQoF+r/77lTNf2ZXQuWx/Kxl1ComuPoQU6zanWwwFblsm
nxlF3fi/CP7mv4yi7kxo5nrtLW++PqVA3Wj+ZdXC9AUwJ/Aptj333aUoNiuJeibYM5J/qEedT28Z
+g/UV93qEr4XvhfT1FzFoyGPq7aqeZZ9Aj7LdNGIIVgIIaez6ti9sVNnL26FFpZ0VSroyCFYbod+
VJLgh2kJ0cFicqHoTKmNKt3jmXa0ib//EQOl2czTIPrGraOQAR6oOeXGN9eRWT/te8s0tNhTEVfI
iOZRSAUFXZKFwoCw5SBL/oKSIjWn2ChiMIJRSxMkwnvEtvcPX1wxTj3IR8phsMIqhZYoWsF46ZhV
Bd8nFtD4hCDdy4RpymG5Nm/51Wsef/5GUTtdvBkhw2tulwcB8r7f5J/3sYXwZtWLQUUae+71Dls6
ooY/Tztj6IPlnsNvoDphhKcajk94xSncDkDRX0AsYVINJxcTR4fsVeBQqnFBHlJaK9q1qObLT84Y
Aih4JFJtTst56zgXqMYJBNaSZrZZcAInLLws+UYfXkSRuZk/RAY3ZnLlTXazPjzcYsj+LRN7zUmd
B4JjMBz82NYYhOgK/KJmGBeqnik5O4GoEL03O5sQ1hTwX/JC6wh3MH/Dl4DutFVbtKSQ7Jr8cf3a
wFi1HUvUmxQ3kw/C3mDz5JUBMdn4h9cx8WAvxxqEOlrFM2vNoK+znrijOv/ABPjrztHVBAJjdoZl
av3cKpMIk1VexSclBhU+nw9pwnA0hf1rPiti+0oxnLHIUsKEIca1y5GnZuEixORmxmqjvUVrd9QE
GRI21op0XmUdw+IvCPQ9FIt5vmICXY7Nvb87+oo+zMOWXuyt4oGAN3Y+4rZZAo2/uBlcCgwFs0vv
03n4POpGMSHDQEC6R51vOqt2F+uKabEqG6VnBauwZGRs7LocoP/rnQbE5NxvPW40qjEz5jPuqsve
KO35jPsuqRB7Ix72IEAH+XxpgZDLRoSo9I5WGJZnGsrAwQVSNwyvDm1j7jHO9Kh2deW6/LKQx5jB
xhpjRweDmoHnWvV2lcg/vl5KKvyWnhzKzyGO8Ic4tjJYL4RxI7JrPe+1O4nm3Dq5SCiQSbuvcGyE
H79mKscZ8M8f4+c5duKHHKHxHP8H+hv9DNpkX+w3r3IAwu+Xq456NLRz5hQ+CvaqPQeY10Wqiqp5
UYsegvbLyds7neKfqU0Xhrxlaa9hNwS/sPyuEZLJ+njdkW7OLhscAFz0LleKn2+0wGakarJ5fMnb
oQmri+7ECItiuB+qmWjWPg+SQLuaeo45JThL3XRPyBViZZKDars/ot8HwpBaoJW1u4vt8TTUPJai
JxlChV/8UWHbPGrcqiA7yAjqaCbSeIrangCY4pL/NiIpGsupg52H6VC9+v37fj760Zj5sdMmpeY3
62BDN5M7V/kTeh/FGplFaL5qN7nHslXxRGtaZSa0HXfY1v0zmHF9V56AsTNT6UUNVCy0hTG0HdSm
+TJ/nCpaBvVm+br+9IDsckL+ujshM+tdJ7o90VWKm7CHcVc1HcxfJqYIwvmJ/xjlDZMjSUWbzbDw
sFsM3Z7gI26CfCDcsgk9P8cblsrGysF6H1bzkuYnDmX6FcySeuJT2xdwAAGhvxVQjj+15+xPyjHc
7GEK0Jo3mlc4YwwAzt8yzJTHGhHWrVZ/+5QmdWQ1o6GAW5QO1d9Y/wUHbFkq14vsaKIXlfC60VLP
P61U0fDSZxDOSughvDjFJrPtgIxCYrSxeR5irqU70uNLHXcKAeBOlpbeb4J41/w7+Co8V+4jlmtE
QcOinkx8RkqDYRzNnTcWIPenO1vTNB2qZFErzdMEBZPrNRbTonXEOnIkDyZqC6djjEqOwws+Awrh
+gT+zq5wvxI5uQyibrOzBYhNXZDCV2Pf0rq5UNQIgh9m90ipODKxwRI+//NiAFwt7lRFNketiGn6
dbOTOoaBElEwjggKWArEAz/JyV++xnjAPF/J1reps3AvBou4hfGRU979rRQCkg1exKhg+wZjUXpH
433lM+cKFRkYOCIN02q+e5N8n95BVBbb5irwDwZt4v8g79uBiB2PGXcecYd126NvYc6FOBDXB/Bv
m31nxrcsgfaRK4GvOkBcDWVrylIotB3AFPFoFHJWrMDWJrH5UfQYlahIrrSONwVWBOpy8Ea9L/XI
ONKYHuam+ASJSKXQCQl5O7NBLAZ6+aosQrvigPWAID7f0C3Qk6tjNiG7BAtBEhXB0Og2IfhLYDEF
zXGrWL4v1/Tys5vUFzSIXcDCKknIc/vpXQIuaeZe4DzIjtq6yUUlbHRiMryFU2uGnUJxOAUnw71A
3F9uWgsGwqOQnvfSyVmirh7YCHKeGzSKQCoA1M6yJRSvwoTp6RWLt88z4/VkZcWKqP/jWsBtaWCF
CQdsUY2zE85jqRTLqFujbuLWV6VaPcSkVXXn7WAi6C8zQqh5s371YcXZJa0STnqj0+gr2TJG91b9
uOrsVQt5fN9CsiNlu6iz0eUw0bqkWdnvcRxJLtx11nkuDFXRy5fbqquwhFvuON5DscxuCACfitLb
PZiFp7XgHxviFwzR/DGBD3JNK3RGKRKE1LIZQC3keTbZ9djALpUbLGNgD8cFwt8POr0U2owLmsPe
94Lc2zNvmNO4/iUsoRETIQiGxQV6iF76XBMsEb7iZnFgYGZK2Po+Uraw0noGiQXWrRRKf6ykRh41
r3v2oE5eGFBpE9ashkcqV6VQE//m7MBpEmXLKOvOHeoSzkFnXDSQs/P7O7TKK02uXvoRLxHsmpgd
fF5BsjBFWuZtCVZnMzGegfTlqDn5d6H+udpb9PdqQVlI/MtTdUGAcmLJM1bcdFLilr1kJHQ2R0Zr
5azAs2/c5b6fSv+rS9WT/t6+LIaocenXCtO87Gu5/XFGh5An8Ei01+I2SHhIS7oeIEdl24VtxkPl
VKAZ7ZN2wM5vkenqXqti15fJeUNg/Yna0GOEb4hA/QWe3buAAjkifL9MfpjaIm99ICuKf8IpTo3Y
5vVLLHrplWCtS0qdBuFHptQHZ2BHTDypeIyyZI6SOx7TF0C98HAFf85arSkAm1MV8a9dlepeKrHX
Y/86qieMUhcWco8Z2PQJ6pZelm1bH2G67fUR8HPliiUXa2nL3y+cwVSrOjztea+nfogKhyTcLR8q
6dJHQp0cpqai2nuEr534PW191Lh6Pv6Ga8RV2lSk3THhVwOxRFP3W2AT5gh38YH9qL94qoZxBchd
qN80IOvitQ7mBl4nZb7yyo72r71jMm2WJ6GAIXOFBDLajpH1N06ghuY5EAvRKbY+GVcJ0yfX4P31
i2Jj+wH0zZZ25yX1Jb1Xsexvy9Q+g/pFjPRuuILxW8nb8fIDTQMD8qUv9vVGa5FcVssvK3ohS++p
L4R+GChbUqjVEoGSVungYyBIeGaypOK7c4l73LHBd6TTe5U7NfOiZ7bMYq81Ishf/+x3Qty/xn4q
9fqVv88DDA4iU18eWkWTlsVPC35TyeqWlMe5azP3ccOt/ygkeX5S8KuFfqPPyYQFT2pHQXl1XRja
QYUwOlZG3q4PlcmDM+/EEOTcgDuPB4FYKw+czds+CY3Rs8vgyb4bWEOCTnu+c7+wetyLjiSj6uu9
I8nPLp5/JzCqGcuxhl16BMZhVcO0OUQED/2FqqGQaImI2+54DZ6OuXp3mPmYk4zw77l0ZqJM/GVz
/eE4FfSSbs/pJU85VOzXsa17GKXdya8Frj0umQ0vs9sudNduT63sGLa3hRBUOoZyg0x675foyifU
kQ+SeiIUFD7Vz36OIw5pUtoUFFCFH56gYuopPiEEpIjLh+Khl/3rUYoCXHhFkFz4ib4teoaRHZMe
7Sw5T4pm9a+3wQYUzLSjtxuXRuVLM332SmgLzi5uDePACF0SwuVCYBCGS6G+ppTyOTCW3VuumeLD
APXSHzzP4v71v3/EZfQwRIDWzlYy/nDoOM2j1sOzmd6EayoD3fwDvkpG2j212vLl3rC4t3hsBllR
na1sY2DVPRIijdPochMYbCfz97AFEqOB9k87NcGeLExfRpaKDovU6g1p5UYQZS23qhXmqR/9JQ0o
DTEt27EFoLbqVQAz+n/L/FNlt2izizDPtkAQ4LLsMCHY5n+Q7d+1Pk4VAABPuD35SHOGFBAdXnCZ
Izgbc9OXqpmEzFsZpWnmlHVieyUr29Wj2M8we3wS/ASRcy1ku1FFVE/ngi/0S9rjEULxocGKlVvo
i599yYcnPoRKvnCIID2o94ngDtpekgm9wV7XuZWDYxixWX3lQby4Y7CmkIvNLK9qLFQ/b2dhlzp/
1sJw+T+adoYdTLbr7ZplMXmSPvjv9xj3mYZoIxtvUOm+3Qi23XEYbz3r5qktX8O64Jxkc/HQgAwH
6RjAE7UHolqcU/4XwXWs+cVwYYjFUJ/c1XZ7xQsHo0ArztMt++gnW1ICHsMHls1hilRXxYyOFNDE
g7oE+wwP6/UGscF42lMXJ43AYn6r1IFgX04xetiZRHL5HOAV+7RRabdINQrHEg2Wb3qHLBwmOCVm
hZaKAo90fQd0/8WM+PzJWV2UNL3XZ+7JlXlDl2j9ogZVOT6kbyXSO9TObjUNAYYpXZV21TEwN97F
VkZkViLQTVGNH2CM1JSTLtQrOGoV3gJa4mXnXWH7SAW0thAg5vdPrL3tFNE/NiqpxrASgO0pGwaE
ghtDUiWBOpHwyS5MRfNW4WNow429QBVb/I8ruzag76OITrarSlXgqrHHtWgPRkVFG/MQl2QteUj6
fWpQ/+R6RmDEnl00kMydDK/1/OBfuEDOrlYCzMVcdMz5ZSbiSkbQfFccPORYABxAjETtAlWX5bGy
T+7yqi5UaS4Xa3afwncbUZavXShGTOqO5uyAPBu50MJqG0ECviZFKvFb1iU5/yQBGh5qqKqFQp2G
SEFXUSTxM1Lm3TFrbDsjV5n7HO/ctcoFN9IXYy2yf5rtS7KmObufKv863U61BWzRByPj7QMxyOXk
fgqu9jYGocH5Oi/8rC1r6CvXUWTIQ/alYxI+IGQp4lg/Bs9M80I+q8pRAvM4InTUa0MNhWjCY3GS
GU23uu601TKm8DixnCpeg/cOjxSvl3xrJS4BcLhl+QkRT4AEXOg6zABt3Yy8ANR+eE6XzfuR5nql
OueBYkeb+hKpy/3StO3z02HMViKHL1TrrV95F3vZ3srzRjyvT3FygXEGjUyjt/ODdQMJ6lC/1RR4
ylsyMZnErTM3A5ZLQXCUJsgVWYkZ2Qpz5TyVFfLqjxs9a6AcHvEUn/z2ZHj1xvMIYbKuMWwmOz6D
V04TuS+kzXqBTUG9NnYx3xX6CT9crybGNKFS/7cS2uzQ92QtRMzcZAwLsu1BnWKCUfZBrdEJKrNq
rvOHVsFc8jTkJpiM26dKchCMsTNSys2lpnWJufG8TAscmo0AZx+8Q5a7n6nXIykSAf+E6Byv1R+M
/jp5IOFiIAbtUU9lPOCIUA9k9yo3StXlzGTGmwnVwz6lGzjkrUB5mX5Gjkhj2jokkCUKOI1/sivc
0QWkKdh6pWnZ58AxA7X/zitfe1cbb79m4x0Gha+KoqyjvqCJ0YItL6Ip+mYdKZgV3NYbgxHTmKeg
4X03XRS4i7iwOCCIZhA2ULWDAgj4FSSkOR1a6wC6m3mJUPWsX9WYtqX2fkveVJRi7IuRdgxIeOC3
oICWwi81Da+6XdCi+kEKxLNy6Q2KL5H0ok+TpeLpWrgkWrebU4lsdW3HCaf/JfMPrKms3jR0c7oJ
5TDY9N3qVjEIq5w05qll8hUbH1wiftVKEtGqBNp7Axj0GPXXLezbMf4WQnNDkL22eKTeWZutze/2
4En7PQI0jP3ePoS1UMe9HjgVHtQhl17103Ut80QXx0To+ZB9vgd/UHMVsBBIHUjY6/Y+KbIqejXA
sL2Ftew4R5TiDhHmqlmEGwc+TU9CzORicvfcXV6WC7vPEqf0vRFo5YyhlOK9YmmbJChTqht/5ChS
ZMz+mQjoU+HEKmItU2iJDlwPkq7Dy8c7fBJd+u4tc2uLqVrS2hw7YGeS1n4HrmAiFZV28B1RmwSG
HW2+/6vo6IiGFR6LD8aagyaFqN4S2MXWA0NMWA1jha6YuGJ9PCXColOxt+ocW8pooCuiiDNcYx4T
uF3+mD+0UMDObaTWBFE2syzCaNlWdDa8QiHl2JRHt4MRitz7XB8/a2TBV8zx297b0GaivEXqbKiR
RgDmO0g6fbc9XvnfmP6XFYYL03sXOoVrIwwHioRtsT344hu5pDI0fQqwJ1k3sAcLeFupfVV9I+yf
OQM6LyNXVfxwLvJsLzAX5IFtqM2R3WJxeS/qCqVMBrldqiacxaKpJoVkNSvocY+9FqDCWbyI8Uhr
REObL48VdaA8sLGJKtR1QwCs0Z3jB4AV1JH3gYRFAQpOjExHeRWwkGJ6CAdpHo5JnL7f/8LRbbGu
C2rMm3+zc08lemx0q1NsfA8OrdxW04hVhTQ8fQgIMjooY8o7POdkSG13zbTuf/OOimoh+VFjWBHe
EKfbTJhQvSHdgXKOZYQNaMtydjCb4nP+f41zEtEtsq7tVftTtoj4JDwmB8dXlG+kLEe0zfZ4Adeu
JBmZTosMyIg3Hl266nrox2qc/Cn3K/GFmXJ8V2FJRcRt5EQ0BgqrCCyZBoCy+E4H3H6OguqvlR6z
xsXokQH/SPJyb75TKZO5yXovrTG/sb3e09QnaZiyAW1sjnRDSkfTkbENEGggaNdpPXUu5M/ppBo5
9szJWQnz1pwhQ4nmIzktbBZPMu2GpaKVHSlas3KQuLwtfl8vViW3clEFF19FTXEEOihuZQwlpb2X
zNJGtpgvm1tV+padC8KusuGZeFUxX/8HfomDDjN0ac/6mnanVzqNtArOJX7avlmWUQRZIrFfMxWS
Z9T6mPlWuCQwouZNFbuBO9lCW3plPtdq/JTqUdeLQ23OoSzR3KnbvpHBvQ68K0ooUL2sMPbGcjk7
fl5neQ20rFwxOeBvQMD30B9jAdxcJl4A/bukQx54b1wE1DTsGfhFzmUWU1OP5qPuFN3+0TgWxep1
265RsP4SAN6HMv4GujFPMxN0moLYQcQr7br09fxFPKH2UXacxbr8Je97JiN56hM9g3ACJSwuvVdt
lyoc9zhQFCK17oqFfS1kN8qJwGt5DpGEGzvTTXn8E/5dIY5fkqxSNPl+o+XgncDbrfUyCo5F3o6v
hMcowGEDn6bXR9R5RkWGgy85ijesXL0K5KnNJFfeL8zFAGBdA0R6GYLLk5kMrDMlXQIBblK2gJIn
ZkUBLFYHAo1R0DhPkIan1ojSruTPwg7U2u78EkB+xcjiHGpLrFsXUYuVCWfXsCAVbggz718gZe+B
R226uDAl/mV5cqUWb7ahienID5H2B7s0y9jbeC1ysH+7XcKg4f3wm+qLc0SIwgIU2P8XXtZG5EXY
d1jZNWerKTs36CmZR3T/OK5jWmERB11L/64dBSYblTX5LdHVlCTlPFL/X2lZA6qQj0rw/YTh2w+N
BAd3mkViWN190wuQ4utDQkhbErqjQYx7aJ9rvU0lPQKO9B+48I1V1OwyP+Z4SMISSMeiiANHjDyA
YKLoDcAqsp+kReku8bxg7YosNJtO1oStnMJpi+v07qwhxyBxi9ocgqlivEQ5bV77dpkxtsHb/vI0
D801oEvFJKTnkbNCsNZCMm3H/S1p+c+CUTjsWHp4BO2H4MSClNf05Gd2vcidupJv7xcaH+ChmBDo
f57ppJmfrO+MXWQP4ky9d8OxLIbPF+kfIRQ+roUf0Sy5RA/bWKpPgF7HFfPdKmkXbDTGOfe6XQe7
aXumUcuGBY/Bdol0a0pPYQ0JaEB+PoUGqrmM8rP6kLN+wfikhtlDwswlfDTSZjLlw+BZIIqzOxnN
649hTMfqD81uGqtBvuHHx3VLND1h0tyMm8LlgGPX3v1jTUQwcJ1FZRYY9UBrihXBm0Y61xv0vAJM
4tOS7sWxT9h34o9FCEFuCPHjHbSvRZApwEbidLnvnFZjrEVNX0FNLCC7BmsKvHFjXJwoJzBLr3XU
5eif6UVDwRNNv6SRPu6giZQw+moEFOTX25ViA+DPKRCDpwzHcBXTOL6biRbRkWjAMT6W+cUsB5Td
dtlppdq59tf0HjHwNareZv99Gu4CG2b+HSsUjLHKQiEDAWLz46kaBER2m1/Agc2RyWMKkCoQyZwh
Fhtxtj7+yHWuObaIbYyL1v3lhA+7GTNPO4PgYcVwRf+XlI5WFwQZgzrphHrtp1zGTucRddQuZi9L
qhomgxzfNNoS1THmq84SBSxfqwB5XOmwAg16DqVEBm3kHEgywIqFLv7yWpbPFhBNyr6MnQG5K2rS
2DVGsNe6Y1qImJi1ZB5GHH73/AqP6VqUl+zgo4BKl4TRI0UiB0TR2jWPNrjNLhH0vge6bJS38gEj
1q8eeyvJgsQeFbpzgca9pOHFiJE2jw3v6hhzVhrAT1cnFSipGGnduZm4B8rbZ4/75xA4s4zk2+q5
cS/KbvKyeama4Qyse8XvYZ4mhvkxiyeZuFYtRFm9MXov5bYUXbVmolZ+psdkA7LfhamBOsivpweV
Tx0DZoJiU7KDOfQJVjx0ZiTXA/yb+Pzd8zswzNO9wUpL25NaxuqTE7yUGERRUY0k9YEOExwGK//8
B4wb1ZduMkcWmnvaqKbhyVghz+A+JqDfwHtzaK8+lo2C3azEqyVEXuGkBnv4E7wqPol7xKQW5KjB
j2mItA2Yqap8n5BoqdV42X3lWjKmvqLYN+4Sg4B8Q4BoUUtDi5aYYWjNZTmls5bIvtqnbT7RuD8+
bswgeezX/CQE+Upp3fK5aUekqWHyv6/NZhbw3ljf01h2ALF8XWnQRkMl1aXHa/Nqnj1+G6R+GKog
jekDtsxcLNpijBsbsq8Hql0+EzKXm37lw1bJipeacF/fR4lxJkVpzvQPVz6khwf6aLlxBKjQMgQw
SBfFkxxAF8jYvL9x59Tx24ZyKhQSWhIYMCcL8q8UWPJePBCPLv6eSwyAQx4Eq3arkjFtgCBmGuHS
0y3f0BaG7PlHL/9YFX3AM2m081TgBCG6OwqYqEKo4anrQePHPDV3NlNDAjAWUoFCm8BD+JumpR+E
upnQk/3NMzdbAQNUMdxkkcjN24EAnTl8Ubc8Uof2YmJkfxB2jITHFKoP84ciZjmH6ITcVoDLbrKG
HpF/idru3q84f5qbnVCFmEhoP+gR3UtJQRdkoqSa78YoDCHWP2EYupTouf7KrMZ9zFrQ66JuBVNN
KuqxN51wcn7OHQtGs4m34+VIcm3hjhLwupYPG/hv7Qq6mSC3q+6cyXoUMC0buB5cxr2BIfdqm3La
lVk6I6o4V6K0nMPTp00v/+XOAk6lLembozzhNg+J/BW2vs9BlVlVz7OaQJF0YvA0nnEspVVq+uyU
s/j/V/wiW4LmJ4VNQQNePJgATa9GsZUXAdczUx5O6PVngifZ3D98BBbmheNA9T5uWUED9B0IorIi
BvAOgloSUIGkVXdB851xOrlnHu7S7VezH0myjr7ym7t3jsGSmaobNUwsOcmhvel/zjowbfcfjCAk
3GtMhlUEyZYNzt6C2JXVLe7/PfiQEhoJHIouC+ppPb6n4Uc2QAaGDyR7HOLQptx74T6oO97VM3b6
ZMs76ccGUm9aWRh63ch0ZxHJKN5l8HxvLFs9Ne9s7yCqoTzz7uYiy9r4D4wyOm05INIGN1aIUtdV
JckV4oLPUYHyFA5U3Mvh0kPqoXx1LqFpwGMi0eOuXPkGqBTDU+luC7OcXuVuOeiRE5BwAL0MCpb7
gUpCHrHAhNYIQvZROPzaqyGqwwHYYruGW1xcKF/8AWgVL8jYD4ecvcU6iTmOxIM/qzEN3ajuuRjn
jTckSM8ieweXhlibkd7EhCNZxyzbjyr+uirfKJa9hjvgW6ZL/NDwLjEn3hyzyh8rK2FfhK1M7dKl
d0WVJFGUf5KQFRVOuyUbVPVuB20AklWBFnwcf6L0QqzgJFqxWoVz0LkRfANgHc3d5CrlvOW65emW
EQsnII4mVlgGt7OO6UjVfM5FEwO4iZxMtZgcF5aLugijC4Qi+3O8f3cqqtELjX3Thtt/GYQoKTGL
EFunvm+LZp23qldyW8O5F5x8BO46PYla0z4B0U9Ed80gnRPq9euLiLRpP/q9UCXDzG6I1bTksoNE
ESXyOXcKMmfIBZxwTmsnVgCmO91apr4MjhsDCxHiYEL4XZ8ZMEUNEvfdo4GpjUUyMRrL8M7spgxV
ALDG5AwuVnXQ2MxhjFnF5DIsEfv3Oygm1OHp8VUcYgtR8oWWhwnp7wcObMtL8uk4EzbIM71h9bfF
xyDZKLo+WgVsk5bSRA+XzvhR0hM7gGlKTTvAPwmG2cO1hyzZraRfY9dldIx4AeB2+pi9h7+M6v7p
Pq+BZO8JUycu+thWB+KKPirD9eCUZ2EOQBKwUll5Mutw+i1qNyHUzPwn1QWeHacfQtHkGpyMlK5n
09p8M7bH4QncgYC5KxwOj+lU/JFMWYZHDv8gMxUbOlxgjiy9UJFbwJDg+WjXlbeFzK1K1UutA5Jm
af+8bNveHx2tRUZgDk1bPy3ZT5D5bCQl6UIGi2pn9DCs/IjgW1/mmNUIFLqr1zMJYhxMzDi+2ixo
KgPmFb9QTwEeTsvLghspDELhkWCt6DO0r3Y6bOXXE1aPX/KeIFn8ffVtcplEK8Uz3f95XS1TQ1r5
5KnTb3R36UzifGavJj00Shav5WYaGe5r/4tsW3USJdEXKcgVGnEQDCgLdPIPs83WCfvAuNQT5rlk
8enksur18BrJd6Epk++mIaZfZT7AmiV/i28X5QJ2OmNXwstjSAHmLg9TNuJbmxSY7/Y7m3UBzVUi
eJBlMc4ZFmUUkB44e1QHj8Daf28g8q1U2RwMPXgZ0Fjq2+DJMC41Z8aBLq+3FsHUoih9x+eTKlZY
lFnchkjyXK8WyukU27g/BeDPElDJBhyzTJEPtaUy2+c71FAC/JZEF/KT1MI4RaqjT5nLNVgBJ4uA
VvSocBgt1bXk5WGnKNuw1AH3N6SDKitxCzaWSWaA3DJjSPA71eIyg+ThNrrZ8k4AiZUyS5sUJOxm
najQGOnRrrYocLJZ2XceDMgjsDay42E5k1yPza18nxGxd7Q/ZhHzJ742lI1e2E9E98OAZIRcpdE0
ZX6G8REgz4cFugWHwMLZirxTFGQwHHX2TnrU4IaicTMFOlZ/qodGE2HCswNTsF7+ifOjIeOlIOc1
7bEC7c69tBM9hM1fUkGvWi4mgbnBn+9X6hj58kBaxMu/Y5ImXYwzRIepSTml87dsZUkO5XO24Z0L
S5C9lcLLnmlJkSF1Stpo6EdSS/y/F8saUvL1PD094V9bN6jm/ZI+RfCoNZ16bEVnBzon7H51NefX
6OErfkIqiNmj/87IZ5V/6tnObZYbeqLC5WiVhIa15DRYXMaRv5UWnTuj0Ync8JQup6vhd2ubdH0G
DTLdjTZpXFpPavyObEqfn/FMmB1qn2Pd+eGl+5KxrqztbC+xFIV1r2Gb9Myug4eHNQduPUtlX303
b8Z+HCMAyUi+4OAzlVxNf+t3dU3VGg6uMkQ2F5oPIyAL6+nqxeYzWXg/22oD/9st3xU99NH9eQre
LquYNrmPbSXzAndCbJ5VT9+fVoe9BkX2sirf0DymWkLGj8gJeyMA5bZhciluGKSbzXx30ruyo0hz
8/FFzzGOcrA/yrmiHD9G59KRcjRCJdcvGJhPU0OXhXzRj4nS6ga1j+541guh+96KfTPR1f0nxv5b
d3YT1TGfR55wpPsl+fTpbYSk9HngDF59GqaurS++OupW4MwH3PwqacnBAqvwMSUxqRsy2lTTN7+i
6NOXOkG3fmLhJd1n23M7tv/bf0czWIK+QklzNuSIS1KeicrkYTx4woghSf0ZVj4MirWc2Adw2fZO
b6M+O3MyVADPkU3d/UmmfFd6N9b81ykQQ+/M3x2Slf6jmyJXfiAsZNgiyNwBKhPhEC7+i/Sxfzhw
dPfAKapQSa4GyhAy3L0wkTb8THi0cNK2jbN+pyubsAzc+cPsdGBVxu3nlYDIaS6pPVYbc/mOOpOf
vD2/odvpr8HGr5m28rM5ZvWzGUnr68hBFJ13vitmIiqnK5cejX0QlusUQlo95CI4GVD4EM/kwhRG
hpPCKqGc0/FzdGH7OEsxbPppGSmA9AeS7UwVpElJ+Xla+vgTGqQoNuXkIhSo90QvQk5uPAkeqmWH
cg7HvjiGYoR8Ywl2rVPcOX1AmJ9oRfdEgt98WjxeLEWKClFHR9EXP+7W704DtFj6x9sxCmf7te/9
R/7G08abgqM7GIPto2+J3zDqz/OHfn0iaPyQxsaWKfpgfpwpnMdu18c6mXRZxAhD2PhFYt2SckTv
QDtwaxB7zlHLs+FJ/ztm5mTwgDUV2J9tiuR6bBU4bfYSWfPwuZY8QnDRXr71CMsCnPOj2rov4ISC
7tm0+I/wJCY4purlJ02m/wI0HIyxngnrbn659zmijro7DJDeBzgor+nJ1hfI/a/9Z7qR5OH47mxj
a1BRJQAqSWpOc/LtVbvxQbSTPNNJq/Y8D6Bi1gWEhAcKnWK1qF+eDmXI0b6PR/lUnLLnqIMtqzT1
Sgku/C60Qe2u/QpiIYjjNjzyXATuYOy9tsWG2+I0pjyAbUCDK4gPCkbk8mtKKOn9WrUu292PHRVG
JI0nka/9g+a3m1SxqNTI2MiLOvMBeEwibidpNnCC7FYk+By7n+UWneEcWZ6jYz49Yc9xENEd7q/y
2Li0EOOIENXirmlyz90M6sgKuRAGLmZU34aT7rwLBXfF7bh4RSKbUOkvlmaDWb0I3BgUinQaAg35
okIcGj1mZEUI9FVm62MfjJn/vGCgvEb/+NffCV87/cng/VKCLCt1sYNP2U5dh+f865WzClN+G3WJ
h5oOqHFSq1GbpTI+vx+kaRL2IlfBZsVmaasaw3w/tmVWuh6A9XA9vdiEfnEFoaDFLc6HvC+akShH
Sna1LaaorqYEPlYX08Xh0YcKtoXQmvaz53ek43YDM8MaJeVwGCn9k/W0L6m1HlC5IOWo3P5OFlYr
ndHw06EIMKMB4IMTyxPycCzzFQVl1adnnvXdeie40iKmKpZ5JTP+fxnMnHd/rBCdAdNbFQ+yanCL
jNX959Bf19cM/Bj+vgu0Be/ZLf8hjjLedbDf8C+QtrWcz5BSPqW5+X9wDzzpcIVGvs8uYqhKrC6/
r+BHNMOKRyKilZsYoCv/Ygy4Yg1m/nPZ9wGjkE7a4SWVThXijEBn71+kgWRcxD6a9sfYiK+lSMo2
2fKO30hmL4KgUmnpGiwWaepVdPBALITfsOJkDRkkebrbqsOcqRC6hYvpXy+L/BTLXz0wHUeA5IwR
xX9aRLCro/o5Hm5cHDnz7txWo7gLTAUdSz7x8db1H0dZ8PFqIyNs7mlxuJjltBF8MtJtPn4MR7kn
Meu7orld0uneBhGqb4X82+6yhf2Z35dOSORDbk0TWr1bF1kBYxJxgSHXhoni0BKgD/qpFEwGrIUZ
xIshZR/tJ0l1fN84CRpBe/I6vOstwoFq2He14S2L4koFT12Tav5k2nH1s/WrbqZVwtBohH3leoPs
Ymp2Csulo0rELabneyzxlLpakiVqFNSlOQ0bb0Kqct7Rw3ziYE1UnwHeheIljQ9fA4R5Fai7sG49
ieUqOTAu+WictlrMeF7we7ZsiGgbjxSCwKlHMQml4o988ONPZL0uenMCOd6dm9iAI8Hh9ebZtJso
VOLYYuVhAVoYNx8NmVar2e1xYC0QkEFoot2/x6lpdIr8no0FMHfhLh5e+rlVfvxQrIdCiHvJD4Bp
YBYBFJc5R5KOwyCUoXSSD/KAlvD3a89qACuTrXoAb3pxzi73hXktef1chepNQmPbPncyyBcsW6wa
4pL5LcKDPTpprmoI7rCV5M4kffc17amG8sALfdTCNa8tcMMpm5rsUqbY8XNt70IfEymViJ+i13JY
AjoltGhX+e2Mr4LDIvmwDZLp14hfE2CY44qr7y8O7YZSSmfOyrv3ITq3pN+FiFD7pGMBiWxeFaqh
HAsWyIA5vZM2VcV2LmLUpA7RamigVaQ2cHPuDvxFJGnxvOeUxglkaBCeTlOwQuzVm7MRELTLtDmb
cEwV+XRf8zzR0WIGOUkP2WC5t6p2b2Q4VSUs5OKfNqsm7GwjfgjOPmJXizxg4zI6DWxP7JzLNlhW
F/1R72WDwZbrMPRheUGyUvaHpmw5C8Qfdrk6fSyjU1ZWDZ5Iw4g5cp5pv9XO6jrWwtYFILWHfdpo
hdz8cGG6oK5YI1AovOCWVlAVqCopjarjjkAkJ53dWh3qHsh4nm+qzFF1xETCYEkep6iNHetlYywq
UZBe5YU+2A+HkbRs9gUz0hmKJohQsLNpapM6IBDWCAEZv/OxUAAtLjLw7M4lzIciRT+Evd6K0u3i
hRCPhEhSLMiSafT4mBWXAUp3lWzPt1v5FdlPgIZwQPO21mweduBufICX3ovAPC0YNNyPqgQ+zqdg
KIyDRxlThovSFCwFqf8iFHS205viWQsoNFnA2750ij/TL33fM4E82U2bNnR69AuOtVA6VRIn53Eo
bbUdlxqQtD3+7gj17aHO3mAerF73h2Hiuswk7tM5WADy3FPhysYKcIXsFCla9rrawlaPbTgAPMsP
aMOtjZ7CrdUi89pzRvTjyL6PumXlLOaJtzbM+f7J16mATzY9WMNy1bu8Xw3LNgt8Hs1XUhQk/dEx
X3SCqS3u0M/r+sR6x926xlDBbDII5U9M6K7p7Oq6LUjRMoM2QbrmDpQhOZ3gyeZcUxcz+tyMjtLf
rIx8tEx18lMOs8JomvdZaJyAsOM2985Y0Cocgr+iNvtEIcrSqSU4Fd7Hfe+Z0USao7fS+XeY7+gZ
isXzGTZm64qobvIGMYVJeP7i7XNGtpN+a3y+4hPBdMJ1Ij1LvZ2vFYbEgZKMAZT+/EmPKp0V0xEs
FYnv/NPrIx2bgdQvCsi4u/7fuJlKjoaxA2mo2vhEduqP60DUIAEh2MgMzYaCT5kbAImHK8QvaDax
jd0bfosAjSpvwJVYQZ3kBZknUBgTYEHpev12YPGQrKTvy8QbaCFrWQR/vJTTM+OH8/5Qxlm1bPj5
fJRFbzB1HEOuziN5DZ8hy0Zoo4DbOsnWMcWGgjXztDB5he7wodho9IzXmMtrP7G65oBKJxZcc//B
dtn+BFCpRe8bc7wpQDZ4ndE6DowOiwsdBMt5hbn2F3Avgir9E3KPLEWbwPluttvXg6lbho4cq3lJ
v7tN643dLL/KXe3xDuFcXiTV2xf8N04KQAoPAK186BOoX9GQxWpmhvg8+Tk6Jm1/KfnVpxnGQqWd
CHA+oJIHlrX/J2nC3kwFtBYzeX8XKQlDkQ4Kc36kh+QutYI164b2i0EYYxPLnXs2bhrLm6ukHB2S
fh3lovRYO6hXYroTLvpAgycsBcEQxFOcLFB4kdZnvFdzLZoSQfvqwjGyaLk47AlID8t2Jmgvcz+Q
gkTMk336MW9FBR8Dvwvc8t0vqbXuoNlIn7Qd/gZLShdd1m/N5Q0Mm6yKwPeQqINoi+RPBdIYyVMu
XcM36R/VRkg5YfVgS2ei7F/BJf9J9rxeJ4tw6hIQFpk3XIkBTh4i5DXy8Y/y7sxYDq/PNEW+2A0U
AqIk1024D+SSwHBP0BXNwybwm9pNPFQ9XKx7aFIKvGXJk0cuzZ09IOuo4QrZLXd1DefNLLpyxhn1
9a81f/Z0ZBYlBZ75qrPLTlQq+jWKYRs75VcCDXT75nBc0iASaqdcjivDYKLmiKFXTIw05beyKl6P
BW8swh4sWRtNWAPASoKbrTcU/juo4y2+fitUxstn53zgG2O0Z+GD8eo8mR1tBS2zwRhgqTI5ugWH
iwPpdoGUC14WvFx9ZkUvkJ7J89h8mzhlEt6TkslNNQnczeyyon7yoCZsT7j0wH7teJ9Ob4jEIFvW
boWc1VoUCe43kgTitsj/OxCv1bIwSKKyXIiCrNaXRRT03fwg52K7r1BW/O6cUnx0isj4OqHOA1Ir
HqZSh+ttefVIKoCLQTDGkwY1rQIUn60oQvLR76tPG2eVT+t/U2mt4RthslBvIilvMZXDITm2FBJE
JfWzsY373K6F2OgI8MFzVjaCVPv2aEaphh8MzfuJuIO680g7ct+mSmBPZkvrmXdJo02BbX4W+pyl
CLUnEq85XiLGVBcxtw5HAPVCF5a9M77m5RJGbRDV1j8J/rCZJgHkxkdsThUM/olb4DHis3fQnio1
qvUNynbOhORT9+UzVcgayEzVvnJOuaJLVBu7nTMdfsPjmuAuzOqN7us62XQbuVj7RBV4p52YkJOe
eAwKd89haUDAtylYR400x/kiQihYuwulWq++zqyJwErq/+6xZ7nrmJovMnKuA7XKr50d5P4wZNZ7
LQI2rr6N31pnrwJoJufc5zD2rQmREArYUtvhMBdX2+Bhz6GxElCi1C1WLynxziuJUK/iOCo6gfSe
7OYyNp4gHIuigJAR5CQ8iOQOMf371VrOVjOXAzO/13jZ03XhoW5Msrz01C4iGwICUgOn0qt0lE7E
pv0x1vLI9+QDYbX+9u1iO98RcauBCapeMoAb2UxSk2DQqql7RGUdl5u6s/i+P8dvq7YvkSwoc3EY
IKWujCTU6owaGLmqdlu0N+jm3uclhIeoZkI9zJGZXoJA0lJTnzrlmGKWkJn66wKkeBK8Esfj3JLE
FxNdyuHW/YIt+l47M1u4Q0twUSQL1qV8ulKdqDloyRzzsE1Rt5QGSJK0cCI8vY3hY9b9e1Thikfi
1gmN3mjhwJow7UWHZuOYIrYn9tvzYXJThKu1g8R7+sAMXw/3pvmKSJ8cUyGgOpJGThLxNKVqCpgD
wuqHLGdQaH2M8BigIyeBispZAYiqr7ItD7rtM0rIBUFKnj2NdU74EsKVeq2ZOnQANdnwiAh6enRa
djjteXhrbNv0mOsRUa0wu6paWOh0ShG9YuHH0i2aBiofn4GYcct7blj8tCx6MjwFUnQAslf22D6b
OIZEuCpuXTVK2f9nLVyVkwPAmoV8ExeVzIUWWwTgip46kZtbYQkpEuNJOKrcCdmS1uQsDrKDfJOa
/OuUL/RAsae3IsOh/AP35X2OcJlYfCQIIQFcHMJWf7Fhqu/4StDFYt3IKWwlch+p/CWUW/QrpFm3
lzHBBd3+kmaiJMR2tJ3C/7n6cVNoTVLbRHya/1LmtGu7miuTk724rEJ5q32Q9ZbJW+H2dh9zuhwb
0lFn07wP89Bb+8XPa9+o6z8PD1Y0hyihe9zHOYZ2EoZ7HyPmpXWMzTx3rAexiQOjw5r5Xr9T441V
H/frR46zBUGQFUTij5EaYq8jVb+aIlE3lrAXvnZhC/b2EJ6Ef086lQtK8n8vLnksr3T0/zNuUQ5s
sVpMRelJXYsBvWBLY9fJLlXm1JWhrYbqTO6dkHzVsoe3sWNIDQJV4y3/LzFgpxAbhwYhheQottDI
w/eLhFoSoPfGogDVSkOxdDPvBfqdOLFNpk5nDHLF+2F8eRWJ6/TKaVkE4GvOIe9g0dYcP9TvAvVL
MzXn7W+I02vOdX85RTwsPsJraeBzD0KDQDU+h/7UgwSariGvk6AmrsLuysF76gJd6Z7nCkbQ5Mp8
yE8i0z9AiR9Z1qVjtaidLVJ5008lBumtlsT9Uj4Mt2nT0vv7JLTKCVxrMT0HPXuqBdpe8KqPtUDy
iMoLldxaKAAleStK8LN5FicHWv7qnKcrzEukAVSsydjdjEPgBaiM8XOtug9fL9bLQNWo9VYx3msn
Q3FVu/FLP57exS+msIhnELNGZVEWbGSkCNKqPESy8MR2R1HYOort5P+Y+SmdcVzw4UHLnxOHhycs
4/LrP33XbSSGgA6/7SjQBZMzYs6YAYYbqJYLYN/6S0ODRaUDMzKmk/Jz5gopaKZlwllYZHZZqIRV
vBel5QQt/gep8T7CjWy/XE399HLWTURN7ywlV0GwMTkuXm/NoDXYk/nxjqhBVub1Eg+bZFNTOJxd
To4etoPP9ZbbXCMz1k+6Zoi46C05jeql0cYyJZCCJc/2Jqb2Raitqyu9fgy9t9IAWOB5Yw1fD9Vn
Jt2+TNCt9omR1kewBRr5to/Z2RC1lVggoQaAcOWitJYt4IFLB//d1nu/4whSmu5zWqlAjlutDRpn
VmMeyeJMObFIEwWYrXNXjIKDfl+lp0ZlH8Iwk3s2ELav7kN0QgkyTuPkyRppWzicJ/t1fCTvMnRb
7W0OKJcvY5dWtev9OYjTv1No3/JqmCUJYQ71/KiyTxeCX7gwgK8hu3LjNfS76SyY0W4wMl1Cwulv
nC3uQqQyV8QHCurq4177jmakGt7l1/CznNVF6Bl5yRrYsSlHvhIUBfJNmc5HzuyHLXk0O7mkFUcH
X7cdUKot+deh1vOBoodT+IykYXSQehp5ds60CAQO1wXZgQIB2Wbbwn2LiS3rTc2LJ6hUgWdHodlJ
Z04feCO65wjd927BI47aqU5CXmimvFt5koWmO0tQaTCpRG9yw9iGnbMQI0AScZ/WQu0VB+Y/vCOs
qJk+eZQVpXUDmQV63jSYevYGaUfc2dhgfXXC/ha9LfFoHIK2PJMEwsFF5HOnFYlGj2IdHuKjoQR3
1RTXFpoNeVSK8gTlAZCbBXajArjolnkFz2k8KbcxZ2CAWV+jxWk+xwcspkc62yP6KnUXR9uL/Yvs
yvfBtTwUJT/xcZeDo62YQhxndJ5GbYScFTXoyVrP2I6XiXXq/hN0u73OjISMPywjVfLu8yVlRj/n
fNJEeWR2g59usnNQuYQtHqwKk67BewTMNc9nOds21e54YWf97yvt2fCDj3C6f17+R1cgdrGj9dt5
arCLofUYtCcwrxv7E80U6PZJGvRWZUDcNodF2u2pfJFsaRvWbezXKocqhUjSWe1DgH+Ku1rfgbFO
WX8GIzYnUMezUIb7keyYK8LyWkffiTEISFexbgTYxrEHS8oT4pNdFFPsMn17oPt7IHMZSS+A8ubL
B45UqRdCRcXVPoo+nY2cXcHV4460qemoS05ulCdX1DjRcBzxgBCyki54d9J5/K1lM1+HoNQwoxaD
m017sRxoWRGf8u8dajuMappnBo5nAbSKJyE29xaNeraQwyAIOZJP7z4RABOGeaWEa5nCizij2DVb
+xyRQwf4MxanIGaZqN+L+3NkSvswmqKzcUHKW7JFbIy84xtksKVN2m8/1Z5QTqSM0ZebwT6qG2jJ
Gb3Z/MbKwRfo9CK+7LChP+GWlpR8+qWZLOOcPWa7xRKhWBE2llJtt1/X6j3EtzPz5vkpBxV+p7PM
atFOc6Ayjp4p8zA18/oT1FTKRC9ouNf/wUB46eGdmAzEtNpWtJ4awQmLD/RE8RFOlhAmqFHzFq7L
waxCMA2ceX/PWB+yOTgoENI6MtifOJAWey7Grz7h/RaHSM+/d7EVGp3ryKYJfzNqeo9iEFYUu8yr
7kagxb2bjYZ5BkkZjInAOo03FZd1hSWPrQMd5uB+tnMjVUbPzXoTuVE1Ef+lT5dt49vIac0wSR3u
Iot3CMB+kWZAmf0Q9+WC0IbZNfo4fpLHNAwtXuRcu9JmTLb6xX+6iJXIQE0XzxJASQ0JOYnDzRUy
dQyieJMZsunyWbsRhKMwbWaJJcZLzYNT+O1UMVntqqHRMCamASupAOS72WgL9hterslEQ8jW3Jnc
f4Hps4/7O9Wi8Q7WDUhh2sLqx8iRNidvNOieXV2x4OKDmLwlVL9Ch4zBv8bxJpXGK3VEDij/l/Bp
s9VnqNjI3FeuXaFHF54aMs9zLLIsgYSgB0V7f5f2kE6X0T/XzTiyS4bSQn8uGR31SBXhdnRX/hlV
ttzczvvCsuqCKIw1iDa2TY4lgF8NtojwvA+ES3WWiP9zUfHCrWAA6AFIc4kholi3sB85r2+1YWJ+
+DXL5k7qu8Be6XBGjsrQjqZqpKvLzDIbgDQefE1mzN0lpC6oMZRmpKTji3XmnRR8lV5Uvj9ZxIxt
YQWniRdb+4LazAyppAlxtze4gN9Xe7iH9Gl1ldUDdzgwC7cntV6vJEIEx7s4qGuPN9UN+A5fyI+9
Vkb3Ry5h8T4t+m06TbEEbgHjDwXkJT1We5UYs9a7OAH2l5Xpz1jVLDrJdalwmMLIL7QR3ZeiaUlz
bYh+xmmH8/cu0FHX9OGkzlpmQsy8g2pOEFLW1+WWIIjnuECAStZJEtZOyoWSUOolUGtSTQ7xZR5i
eMdtVT/qJGQ7VAEZeVtGvJXLVDIM9j2Q3JYkdWax6BOJRN9J/8NZSN/5ie0uHksE2qASlY8AZxRT
4wwjBX3EpmIGB5Vsol6DbhqZpzskJo2YAhRqmBtJ2m1gPe7KqZiYvTTJFOa02VKxsIHYf2C2ySRm
1SsGSCKU2CBKGS++6ATYoOhP2PZUe3mlzostftX+syH7obgNsVu/cJXSibIC+RGFl1YLlItCoN45
Df6jjs2fYwTY3GN5n6YFbbA+NWrCiIsO3x3p2vYsomZmFYRHyontKYMfYktgL/hX96+ZdRX8Oey6
BWoqlPyiLjZ07yIxCfjNbAVFlRaGW4/IEl/3y1Xdmt5pMRmrY+KWgKmsMSBP/D1XzlFn4xQX22DV
yj4kEYjI2s5k6rLj+v91CmtEq+isLoVkI3sGqlJUoWKbofM2mCxM2NbwQ1UBR7klNB5Yc5cRdErc
8SuUcMQLCSdmyBUslnFxMdVsygHyNuDObnEw7tZABFw6tXMLNrqrMn1m5ExvWf06eit/AFHhmsvf
hVfnR2KPQLQ0KdmZRtT3S1Ay/4A1cll9XlIdt1FCSXZ6uAY6L7ppqg68gUNTs8dYtojD3ceUnotq
LFL6c+lnK16lPBebWdbdQEFJrVQbZFVuDki0LJdoE5/tXfmRu3VtEhiyjGeB316bHLP0kx91y3ab
9on4Mv2GeT0Q4wvI7/KuI4SwjxI+1CKxAwP0YnwuO1EJSHqqdly0ne+L17YIm/nbePXYjntzM6g9
xM9fnb9XI+FRZ2CM+HUQQYzgDYEOpEUFezoku3yDjNDFFQlPt15nDW3EqCXYe2GRQt0yIylFnrlJ
t1jypQUVShbzw9MJ+7ABZkojnKv+RU44CHcmH3QO6XBRDSr2XDj/fZuFJMkWQ1JfDtvalSuJ4EaG
HYlrfT3OZVpMqBaZHnzx6/KZGN/0ihdYF9fFr3OqQ9maInGZZmGBp0T5JhtosvAmi/YhgzmLAL8j
fstA/he225AezcyQ+hm/1nRUyoIGltflXoWl4Hlz5orgJ4w7X2i0zX4AZpkglAHK3hLR6psByK+Q
o2myxvNv3IKgjPE6RJmNKFxS5jARX9iM2a/5Jp8hkt4EZnkxBD8JLxrBpBzN2rsyTvCzGGqNTuB3
WXI9DNEbK7wWLgkqQg2ga9VEsBniJfrOIiCKlKgMDLUFK0y32BSxU9J0/lASZisIWAnYqIftkRYj
tm+ozz4QfW2q8kFzBqs5V0VhSmRbKhS1EjTZqq+avlmDO4o6U6xQpdIORxeuC9+y2u6fvis/DrLN
858dI7DZGAXY3S56PWePgaMCOCEYcEGYOVbvR8SL/uZBwqLXt9Z3qI2hi0Xi4ZE1bHWHAvOmKY76
aJ33gRZj3DOw6Cel97FaghpzlVHcNNH/T+SU5mAixoXm3p36aowuxk0lYMoF3mfOpRbAlSDlCl9D
XLtgdf5KCQr4Gv/73bchQOVnoFTGhCaSpyj2LVvpNU6SxDrou7J2DLXVIJynkOPWUvrsZW8/AXjV
8ugWPdEWEXcFGKjmbyUzKArIqsPvj6aBMZfbj/PERkSrdGHy9XKEdQ1/ZqN1xOsGD1EX7Wos8/BV
i+19SjZ+ATivQGNebNEpWyVBVl0BbWxyk/eMWPEH1YlW0u5Z9mqfk4Yq3EDV/Iw9/m4jC7qR3+xr
O+aynj9bpW8cmgL+rtX2YLryosnTki18jmox62Z6HThFTecDceQOKaTtj4Oetm38aieFjS3uivUd
mmys5tH37ImZx9CMTzgxb1ydktfWu0pDkQoc2LZVEf/o3qWA4L4xgdfHViaWY14dwsgam/+rvwqK
yuaLINJ7Y4Z4pqWTdbB45MKnT/rITpqfFeHkKkxpXcSPfRLf0IuasTvIJEboM+3U1nOnXklieNjW
nMKOIXgUpokgRMQ2dgkUek+ch4ff3QFPLuu2H9Lsn/N5Am/F42Rs1Xex93ob8kCtKMQwW1AAJVfI
O3WERz0KG+kO+xyAkHL69cFgpMo9+RJAnepkVdMwaNmNNSMe9wDE4Ie+EURVEnfloMptvAP9vOgU
DKPC8kmNrOW0n3rmf/0F0G+B/xT7+6HKtssmWyNlHGDA1wh1V4uacruq2DkS2ajhtImumjJxSZkG
/gDoNRorgnomfXHKFRO1nVBFPW8diJlboBfqYQ0U8vkNDk55Znl14mHdgjzrE8S7OSVmoqRz9yrc
4S2HfWAtHNWoiTqz6sA2eYgdOWJdWSJwoeaJSgUx5sW7HKYVAWasZqpvpCi9k9jqv3zqqmMiqtbc
I+yTRqXHRGRfGu9K2q/vKbFv0hNBURAenIdB09fUXq2RKLfWZ8QZSCmXMPX7XriZA0gbPghNg23e
Is47TmrGj3cBUzJrlj8ALrRjfRKiibsKvAnKB4m+sRM/m7+f+waYoyiGevy8mwAbxpCTHUsD+R2B
oWRiHm5WF009JlQLqfXpcfIWkb40NEpEJOAo9rFHY5drIoO4fzJYZVrNTzTHPMPAIsSxC8rXczXX
cfXTaRyDkYlvyOuxj44Z4lvyMohANSAoQE8f8MTLwA/XKWP0qHhE6aCdVH2+icEPJZjf8JJjNIOR
yeB5OkivgevfVuB/6le5ZEZHCP8uS0S2U037HL8WcteURM0cetBPJ44jIr7UHPZ7ZXdKVvuM4+xh
hWqIf51PRtf4tO+u+29yvXrtMLXE42oYFuRfP0mtPcKEcxsUajQmxbMU4ElL/lvcuPmYa06Zx+c9
U4wNMiSkgYaWCKRmHVaIp1vVu+/FLmol3PQw+AykliQHbxiCQ1zFgmMEe68gV2JZhBB1rtBONSrQ
bnDpo1hhB0kQ0yiDfW0AxZsYmxex5uSGXrs8+qr7y7+VmAkae//rCCVgJouwmZyV9ysYmZIioKAk
Wy5e83UqPsr5DDAVGYyy/pbcWB46/6hTNyU6j5QwB+EbXKHBDfw1BPRWdBXDCehplEZ+tk5IihNs
ak+190UU5a5SLbILrF8gJDIa1Iws/NGDGrat3lqsXYNJCmIJQZK8nQWV2uQlj2/BTaZspmcfo6BF
FBWkGb6kcRGvh9+ZpGiF4Hu0PpvTqeTwHDSnsg1XW2znMA0kLo02VXVA/lfSWTMb+15nGGlgYHbM
L2ho7Dp6J2RMLCCJLzUAQKJi36T/G7HLCW8ogPhwp4tXCvx38SUlK7HXEjC5TUTnBTwKf/CMHLTf
u26Ncy6Ekru3jIbfCyu8ZEYAyvRCB0GRojUNXP1o3g4kFtPIYi2+NV9sHT4qVfg02siHGNPExemH
9pf8S78bVJuoHnTOblG8EGpDj4irAE7ShG3CJKxWgpHs/uwqo3lFvPXBFZL5mxpk6TGq/z0JmCDf
2JTEhZHKUo2PtMRd1Lr8jkBf6iKfxuOo8sKPOI9hSU+fEpfEhTeYTRUGcyXW4iGETFCrmn7Dt9/y
UMW0YnLqV5OOvTqCHujcFG8pLY9bl5ON+8cIqL7fZlzT7ah6tzaKRIKR6JvJlgt1Ql0Z7qFFj/xN
kIvKYV4B17Ejy6AxdWtOm5OnOKnQOj0pmUYgsObg4IFhC0KKjTJvBm88TfU9O9je9OyuvYI3Xrp1
IxQIkDIUResmG0BbTQdi1wBUq2wiSCZYT6IqRSGkIr2Mm322aLeBhxZMoyuXrOjUCfLhxJOd9nmh
F1Gyru3vFhnG6+oIiDdosXQYUWmDlwBC+GhECs425nhLrdRt1MgBc9fWiCbqlP13UpQCiQgcIFDp
AmG5SdafnKUA0cOwMtmE7OpwkswYCo5RCljt/7/FvMgoRE0EBL9j1WrL8qhcuLb5Bn+/WDw4g5y0
G/brryUwUf1nwhdOfxn7HSnOeZrlmOGniX9MShetA43URejQ19dKsgRiHJC3cGorCCIdSytTH0s3
pmZkZzXSoUrSJLPeVCj27QVtttIjK5ouNf6wJYVsctK1EoFelhZR48e6o3LJHSw/XQmw0TRJxhwN
ccmmEAwtr4wX9Vljy/bwjXlfD6QxpA1YImoYolLqNoH6JyIFwE76dzYljo5VRvogTs8pUwohLD8G
khDE32XqT2GnIMw/BqNH5qPlVWU6sJtpeJMl9hIQaU+MjAJM2O5qhwQQsvJODROpAK9ewfDKkZkx
wG3yqrhA8bTcmLEvQwLJbkll68VrHkxz8Cce50y6vEW2/Krm7yES+NWJEpVf8cAmmiyt+itZ2kPA
QlEotLl8fUi74qVk3FJYhHK58zWdFHR+c2HlGR8148bNFyh0aPa3gAjf4rXm9H3Tm2QjFXr8mbSh
G+0E3yxO0FDWyKaDKmM3atESoZFXxaW08/7/50pKoDvn2wY8/IQVNhZ4p+4jijB5+gmmCkf1wiS7
CW54QgN+6QIKNOIBIRIucXoxqQkmHWRi9P0FMLzb9228cIwReMXvkGL7Vv5pC85A0pq27EGca3sA
lGI37Ilkh818/uvB9JWbsBfCGBrbGm4dc3Ae8f7S1pC+u0BOBzad5MIy2NCd415p/0issgjRWwSD
7I5SRRhzL7e100mjVqMjJxRfmatyZhnFQAkl2hqnFmwYUHNhtefKI1ZMUsfNMVRdrq5vQUwcN+zT
f1BWb3dF8jvycjyYq9vOZ4WfI8u8lv7tdzJpl6wOuOi4iMh4icgVTqjySxelb+akYT0BiLKtZ3jU
8PmWn9kR1VKZzUUM+BCWwZoR7jAHaIZJB3oFQiQbkFtnxc4i7l/DeMmtjwdwSexyG9VQr3rRior/
ELhuS+yoR2F7JaqezwGqmu0hdlKbdZ1xJiGVbc0eN7Qx/3Es3VylPyvCuIBk2kXJxr3UOmMsFFFM
orxt2lAQhQh0IIyl9IZtgpaq9TywHF9V7x4CGRkIRhns0Yvq1hq3OrFLIWCvuFNWCK157B1kurQH
YYI9fEetoe0T5WJYHIHuWLFXbvkY6UWv/qhkLp0MpRC5AF8Geet42Xuv4FuMwXNH23KbnfHiwNKb
KrvKiyRZcRATkwdyx9KuRnV05l3lyKbtsQZQOMRHRbdETbQh/D+degVTjsr+C8Pf0e0tioBCuF55
OOIg94Gh6BuCkSUEiwiPKH+PVTql1HE0iyu0+kie+yNG/pF8DCmzry4vVovDYra/YY7nu2emwLE7
m1WZ0Q8Yb8CmIIbWGk74D0B4fJG5ilLAYWWwSeYAmhVz5MDUGELwLXIyuxTV5x1f3iIFMfl8Y66H
tM/bZfPb/Wfa+qNqm2PezIIh3DqI4/QZlt00os7X6nyrWGUI/7Tf1JTQKCmhwGURklxumPCLgCfs
wgsxgGRPu6wm2XOWqCRWcJmE/x1p+kFqZEuCD0Ph9N8aR40PncSr1JEa5Dl0VNZW3HdKug3UFWud
RPjNtvUFeoudL8T5Y4qwj7CTQiYHIIoLILCN3sXF0WgUfweJ3VOd48ZuZjxMaeqfE4VmKpYuG/1h
3jbIqv5W3WOFro2x4dVqS4rdrQ5hU4ZD92ewrX013pOoMDPhVvbwO6wEODwEllofHBj9Yfp/xt4I
kLx0MlPXScxLQ2XBhA0etRCZl7MhZAZh9YSmS/MXVp1UIfNmc8/PI6qgMentTSY1+MeEtoGKgFdD
id4gllvvDD4F2Nm1sQkL7mMfZv7KUNnPt7OdNg0g/wA7wxS2Yqa6RzV/HhU+dn/mLMDjlLBhJR3Z
AFuF6YZzrQYFh3OCG4ErURyOPPQgsK2GDMj0DUYajboPZn12rcpvjEQ8SPQ8sMVqy7ZSoANATT6O
sNHioPIfK56NmZpsVyk/uKcY8JAdzQ/KZ5UUrwuC7Vlmsdtoi2vIxH5Uev3wwLUNpmfOhCZz2B+M
IYBLg82Zv4bI8ZSAuyEjw+fTNi7AYpPQgc61TY1hj+tBdixhbaLawS/56suO7gEwh6mY64gCOFPj
ye4KYqdnBCM4D/7GX0Am+Xckq3kItgOkEKmAzOoj2Y+ea1HcM8te6Ci0uimwJ2S9rwqe92MvB8aL
GLX0V1JbALJqWV9txbIGtOKTct5KtwyTx7tyC4untXbSJUfZFule2+khmbiapsjD+P4Mop/y063n
DQOU3W0TTgjZmZHbIiJ5KLsc8XWBYeN40NtJLmlZGjTOCp/IBzzxv2vgm/8OE4f7c5s+AEOQoXAF
IUU8pGMx/VFi8XSUP03RaB4J8umfptZ0qt7xGHjiuFcymJxv3gxBKHtYPHpr5+4LOgxRMi65Uh50
ys1S2ZHWZTJliYFAJvuu/Gb4U5HnIEBtDvm46RaqxIt5AGHxKhuB31GJhnKkx1kt0dh9yl63Td4O
MkyZn6igQcwWFpTSlQQ8LrjHaV/TvNB1LeNSiK6fq6R7BUTTs9aphHNkRhTsqCnjQUPgw1kTYb2u
BNf3F7LMyfyc5PPV96Xpog9okRmpqSj88pZDqXRazMH2dw2Gxtup0azLihY7jBoBoxb1UC61NfiS
Ad1dgmT2LXmZ7YLCHVpaAu5yrj2YT7HC5rtQH9gsQ3HClCuHYbOgijqPdzjFSDxHorPbDjFadKXr
qvJkoDg1SxiGsb0lUfcN5uDUxuYjgR8M0zuICu6EDXLZpDyGrEggrn0CPlMb6WtU+jIlG8N332Jt
1MVc8hiJEaGFf69VxUOxILaimbRRmoA8ft/lBVLJ0B0ERX25zOEA46Qow9zESIsx5za/bQn3E3I6
vq1KY5yZxd8CgvOF7fxW3C88p8j3Wa7ZoKHwhpWl5W8EKrVz32607yx/ud+um7qfwMJEa7/jwd9x
VrrKbkWUtyo103rZcWgPP3O2o4bJFChnpVnar23GVcvj2JqAKy3nPObemBUIN6NWE5DkU2q/vYT2
7DyotrvrWzJT6kXnYNW/M3J0pM+qx2dOq7Z8NGfzJ2Bx1Mqg+ahLt4EcqhWotzzjHX6AXHJ0xgNx
26KrP3m6KbBeSBKAEEPd+r2131hlsZPAFVX8O0KCtFz/YzJbx/J7q2H4Kp61r7N7SafZX/4XB4Dt
yxfUhqAE+vZgcWy7KB+oAnpOlVLSBaDEoXynTWB4Z2cYwInOT4gM3Zvqq1f/bwT22bLjTGY6AZMW
ZTSKAMBy0n7x+r89r3bZOXDAqzOfGs3NWuywI7KACAr7xZF70JjHNYJ7nVs9jVcdxUMokQsG+eY+
CrAUOGBPa7OYQBAig7CY10nbNI4Vr4p3XALKxifX+bhIrkMCLmMRUNpj5ZWY0j+/XDFvDe6DxtjW
0s6pCdmL0IP4ZR5BB87lop687GrDnDiWZF90kNl3+xSFBjsnmPgbE6cqLpFjb/9vBumi/arP2cn0
ezlSMQeBDIl3wgkXMhgARL2MIDwsQ2oktijD5px78nzNltZohN1F/omgXmTFmfzL+KJ03M9FPj8K
UMQCuermhggC7B41FUa8v7B8y1I/azBtGEEMjlu3Xm/wSkOp9vmub1CnEN11a5sJt0jt5ywEHlDy
yHJN21LgKd4s+zeS+wDD9w12J07NIExhTyu9T6fEZFssBSwcXLcku7f6APPvCAxW5NxM+sDjVmOT
Pc4Kqm39mSEWhgoqf+EpCZku4agEFeeMCaN5S9hppJdchaTOslh/VmLZU+UDkKGhfm3GqRPKt2BF
hZu3HLkbzeKntRr1qB5Au6ORupYsU/pz9IcJ7NnoTHsznhF/TQQCBjlTSXtGKNhNgwKOjnY4we1r
NOqkJPt+jvbzH9HD2ACbIfvRT4C9NslyppCvJINpNR7wzF/oQLcliYK3s1Aurb3b8ALkx43Nv4ti
lEqih0Wt/YQd9ySdOmMd8iAuBls/TGqyOAuUpJS1iV6urJRV3uLguFgeG+QM0kkZqXsvEumOo2/u
Nk2CLA5kT8gV5RqFvpy30GF337CwhxKrGldBuQUjbEqsI/hvcpSoWqB68RL/bpwXyTCxhKVFnW9g
L8wAKYc9LLyl40/d3+NtJH9OqW3s2zjyOHv3pRlUtRmXHoNW1e3N1EX5ROriFYuZQHpUiQsCytvT
8y6Rw8r8uyeKppihcQ5DgO0ltrVAHgo0fqA0+m6HGglVrTKE+m3JFcSXUvxLJnRhlz9APmmrGdvn
7ZHh731WS45s7fc6+TMow6GOcq2Lc3jJak/jlWcixPxXuP45HcMSDLRZvgZUBRqzL2fo+Qu6ER70
upa+kEDpKsX3Hm2gnqPvZeKqJwehk4uwnaoMvMIRi88uMSadVqfv3rWs4tmkEe8VmDIAGbSQ17wn
1RjsaJ5Kt/IV1kHW2SUQgOJWMcVtYKClbTWLSY5sCtQyapQaXC3NpOERHscQI3PgzFr5ad2KOlzo
Iayo4p+du6QUHR1lnb+hTeRqq/hnlBbLHajgg+3PPbB8PsYDHoh7+iUtjMjAHNYXwK3tTAnIbGu1
2xy+Ep4ghsiwxRTCHwVd+toVWS4LF6SYReMCBGyRnhNeo2UiO8Nq40NwLc35fJdmIohLCfOoBHph
k8daagKrcO/HvRyLJfSRx+CUlZ2i9nH4ms4zi0mtRiatc/DuTp2JHgoCzgd7bp/P1T2z7+SEiU2+
lkiNN+EMvn12U+yMPkIzwLaQ0BFHCEkY6ckxUixVcCUlTIxcWoYeSvWPndNJ6sf6gE8Hg05tPWSM
CjYN6vlzJ9NIfMYs+20jzqLqE+YYgDxnEsHAF8N5R/8oNAxTtra43ElG06tkysVUbpLAqZzoyte6
n3uB3AH139HK2fw/PXugqXJa4dp43GEPtUBS5DgcZ1kDsr0vmVWr7+9Av0kKXokIVjEWGN9V55OD
v17zS/86S+zzl5Xq6gOGkHC7Smw+qgH+dYZVlWzL2wszURHPi2S/dUQgW60T285W/6W+O9ZM/vH/
IA3klxpocepxDGtRxd802ZhLDTsl/klLo0gkJZYBYluYJarclMectbRhEM6FTTJ3whIQ13kQtamu
dKn5pnYoFzZ+/AelVpC1VkBBmijiNNpgNb6p+MvBBuK7CdXvzMGIsspqlvSn1US8/DiPZlzGo+J9
uowiNllVbD0/7DQrMynXIATirBJeA2WrNpIECTU4HEOgeCuNqX31tsWg+V9kii6argQ4KTbGs2OG
DOTfaCWM6EeQOM8uxWwS6ddGRF17kQ2R9NNsVa3N9SNE/0Q81QS3nVR8i659ODXku7q07xk3QA96
3fVPC7Na+dIEUdpRxfo4bLzbjzqlOVVJqUlsSH2ZERff2ocHwWpE1AMx7Li0pe0MJxkTqYAb+0Oz
ODZ5d0utA7jZ4Dpp6UiCG3IkNvGoL2hRzWPUZderbwjCVjqHu8i33RNi4fHyr5UK1uzvhxdh1ga5
7hkMXum7F6MqKATc4eyoyyxsLLq9mBHQWaBmPU0vXzXg48RSFo9xnnWe7VDplWLZgjEwMAFxhdYt
91/a/Ya+cOBUXVBzZRe1OiCmBK7RtpamLl6aAFVwpd3CW0nRvgnmaHaXNuLvXlyiLGjNzd+GFjs7
y4Asts1VSIjg1lbLkjM1vowBre3KawOLN64LLJ/7SftSq8N+b7JU/urQV73JBEJpk3Y/wkzULBmC
TXfaLHsORvs4wIE+a5XsxbsStel1elXtDh0aMccaK0re4rriULnK2hclLxkOyaYr7hwkE2jqKEY7
lUCLOOI3TzxWQEkwKLI+El9w6ah6+OR5ZIgDjWXQGM0hzT07ji2EqJqTAXGM6YNQkXjJQ8AsAG0+
o8VXyuKo4uFOUB3MhQKcixzAwdsZKtzdpDGUtU2X2PdEVMH/14oq/TAP6dYLm4zj5Ti0uumnjudy
MwfA29qhvnsv02xILZE317OYr0tfMY3GWGcBGKyoWxPUBF2kCvwxlMz6B0e+x0x/gS70VK7RKUOc
Re9MrLuBpUCCtmqA1T2pnwt6EOe6oaolDpkW8wq7bYGRQidwB8QHFtI4NhkDS6P4xPYRrEcNsY6h
P/djAMZS7QD4T2WVhVR6+M2ZOx0rJHjtFdcK//6e3P/vV2ru9oMAfsmvj3mu0Tw546BJOnKa7E50
jPa6F6nxRH+JZ0zPGugxSiHpJcqOiWG1Q7IjwmwK9nt50Yq6R7tRXlPph+WB+OJ1AJgAx68IrohD
lLjWe1YHdp0KdKNS1cVE6vwuqIZ6MtiWbGmn164zFLufGL+EpUblPvzdYqv339uSfz0hIZsDf5+V
8kYa0z89KWIxdhgY7By3KoTYGiFdEvx78BpbUYljH8J61gDuLewdMWzZ37NfkbDekXKaySUzAb8d
Bsx3OA6QhIyncY6GcEz6bWyt/XJuha6QY62dJ6xYgZ3ExqVHOX2OzI8loAsh0RUP6KWu+3nrRJwL
p9hiwkpqFi3k+Gottwg9RmWk3jiYLcdTMj3i4bzmmMZcwQNLEyCEEkNVhjjGZeuGEzIADeMDGT+K
hxeHgqXt3qJ9r2VNPU4FTfJmHuo8U0fjdXYjjwnoJvmYYmTHFrwp/oSinUZ8ihRrXtjB3v8nd0bP
75hBO5worhNjA3StJYCs7BQZcQ7fRcFvnbBiVl+CTplhi8sZofjtOsO5DluP8z3S2BDYkZvP+d/p
WvWiVrcrMCHUscSw6BG/YyjevqF5wMpkQvymJhP57KZMOBlq+15bhgDTauGmtT5QrKShwFcBwv1Z
PKxBN1+PGKovjcBjyNf7zaMxJtd/gsfcyaZeQMN9gWMXNHzekpc4Th1v4ls+CyNexM4LYb3lgwrU
Htx/CAb2hhUgbuQy1z8Ex5jz1h/56q4EEgGFPlM7k2tcFuI9HCVQH14dX9ups7yuzqXayIe6h9/F
p67lBiXUzSx1bRLhP1/ddwQaONSkeW5/kCPBRJRbnZytzvl7nH57w/Zz82kjG1LCd1Q4aGmLKIqk
JxGWramqxwtEQnDYrrQDufYXEKREfds7rgfyGtR/ndWD0QP1fQG7jloTcRoJiaLSeZBc0VTeFsmB
JOYgLhE0BcOl1fwEcz4CZYIyGdil1Bo1e4h9Oqj5Z/U9Wd0un2CXdGZ8MAmZWgv70tuPmHkXzZZV
xSdZqNdJpYTlJwMaRbbIU4UCLLmGFZbSxe0LSa7NNUsjYo/QZBTthK/YPelvFRhBtHMccg/IKmCJ
YyoDZR3vkP6kTaafcMYeleJ1EranNyfptd8XW5VhDhVzp7Fd5RSJJbTx5ioQeKbGJhYf7phXPTQN
I/TYe6EXFGDLnOGDQmitzhqzxViazSG4d7aEZ/8vfNdDGxnU9kyJQhk9LV8/LOb3BFdeJ0dgflzr
PmbcXQUOT5DCLbX9S/1wwYDaW1suctV9hwA5xzNlsk+pXrjp6+IHpjg2F/YVA88moTOilMiBW1F6
YuTH/IDNBM2jwTyeWKo7Bucz6vBMroEm9tlJTC3jUBJTYAsiv/YIb03k8tUwaHAkDckTz3+c4lL0
TOfyVbGStA8NCmsgPoDlDphHyVr6WRev1D9ddHDG9uimAh1fHGQekkiiJTs9X5l5nZcvovqwcvFa
KGwSDi37LbciTfoJdgXZVPIhi5ALVrWq9EZd5xvhnYmClxOMhh0L9dGaVp5aLx+WGgrVJnAmEI45
MRmqSaWYMMjHOi1LaVwYWbSBLyakbvB3OdAmSNucA6r2IloFqSWVQHAnPzfYQg+AYP8mAS2CViip
3AwdQaGE6CJRGgPKTariaBzcLU3bYtZ4zSRhRIfsftRIcUddUk9Pyh8nNDOE34ZSNLxHZdCO6iaH
LxwLiaIOAFbqonAKLdBMFXhKFbh75/o1T+7BBV/I1GOPPeXqsLaiojITu02wueJ4dP4rAZF2hDYe
NDSsfITNtAlX54Ah90SIMY0s3eIPdsfmEbCNEfTnDJa6ww/y+HCz+iqTW3B6PFOLhKctKAB7MGMH
1P6lHYnhuzDmE5wW7mUnGlVzSevzmw9G/f6LYJA3nCiJYFqLinZ6MjwJ3UmauEGeFGHB16T/uhjg
4wuSUwHVpAj0YyoyCRJeeqev5cu6SPLk7ysKMzDpqlGcoIJ5z6vFhiNTTxh7/WGJ67MpQ8gbg5ap
ObXRbuI+tVwciFHwyWJL8bY/mtECYcqnRZq5R9ApREQ4c490Qaxa45VMHtvS0JQlZchTIxZaFjBg
Ak0bmr458OwtZVOmq7J39Li/Iy89xeKx1q2OOEfxLCME7TvxdSGI11P1otiGebUQj6XRqRkalWPc
k9Q0FcXEX6+rzdTtxoSMt/cYjS1PzLMT1BbQdHSdStgywI7PXHSnfZRXogK4BjPN2Y65+fpEBvw/
tW0HBsPjpW7IKfQItxFi1bZN0l9JsVFTGTajD62RTZg9dQhBp0QIVCZmGhtax8EaRhd6bG5JjRHJ
jIDNzWYm989C6jAkzAV63nDsoifS3p0Tip14iOrVPclcRjKkA61ZbzqupB6kZuHEz3TUq/Rxi6I6
dglhrKl3XaqQJoezQ0OlBne+I5cg/et+9ThIFTmqjpx/64H1zvoz/o46S8hxih5bMhUxoC2uqGAu
MPiRE27OIUmBDNdGODbFh6ewrdA8NKKRk51Jb0Idtu9KGaakgRrCyonjpTjvVSJ+6e4wqSn8xe+o
khEnMtFev/xsy+7tXMTgXi8iwzCzapWGGeMwCF6EvQb+bFZ0hhQFYHdYCxAdtcAJBsHY5P8JBcZ1
MgWc87Yrwrq+E9VyUhpyQwpyUFFXpEkp24mQZWJ0vdZB+g/ZPeuGgk/yS9o9k+LbHEJPjSipwd4i
oyZEhM6wXt4kbcHi5E/BhvVpBzzx8xl/1JmpYTHpCk+T6sv38gk5UN3Vq58hQtNYWozZriR8GJGR
zvJnSFtPqLSgcizjAWdqrl1FBQ1PM8S7mXzrYYT/ofEmUo0Q4ua6O2ujWl+wgfSIUXwIjKTWzniO
urBcjZzKak2xIuDJuY4+ct8nYFDFMO5LS6cx25Nav2JJKIGgeu2zLAtd2IPtUxihEKpDOvYVt0MK
1ZLcGXf0+YRA1JzhkpdsgnoD7tQEUxSJEOzafIzm0D1j/DBZMimtRftQM5/RTxsyNcPTFcbmrf8L
PvmZTCvVXL8iIPivehIoxjk4CYr5ulquzAfk1K53N1WKEq7OsDXwWQqujcWrpI07uo6RrPoYhJHV
pKbwdihMub10TY/dvPXYUKGJh+Xui+++lfwTZWRB/gMryUIYaqzQ28MO9iGaiCaR5/GlgThTFQxe
By5WtQ7uBEIYVfe9dLFAL5RqCiNu1un8tvxuspFhjGnWW0JWWqpBuIi2JXFGtLWieJCNKZbNQoy0
5qcuPgKddDa2DVRFE8QfkrpYKiMHzIvwkoBoS6IHUEEjnIYYbgHum9ftthQWgB9m45eBMNR5a4KX
rbSaw5xOTdoQmsogqob4OoxfUB5kM76WA962y2g+ovg19vUR0VlxbGHQeE3Y8Q29M5qUktjR+lRD
sZ/P8PwN1wopdCtYZNOoNwQxnX+7ZB5k88V9Xm5GwATrvuk5zUuStpP9IkaOv8aTgqLaZ7y87Rv+
p+qhoG65e3MzLb7sBDbAxpyyTmOiv6oZAlC+wMwQKDSa/ydqLXXDdqHbE04Sa0h9RiZbi+Zxqr6H
yrscoLdtl2ACpvByPCI0A5N276e9rZLh5LKFC0r7x0urX6O9CIO/ym5OJ29kUmgahlCIkednDY7I
3wAkMIcvQSzlqeeDoUoxybXghg/xuP915SJ7lWoQMPxXZhQKFsiRrUMnjH6YwDiot4Zmx81HNDJe
ty9K3DOwvM9sPcWL0CzAEFV3I6dgxECrL5ThvFdD++t+T09TK16fWOK5b6ogRPj/qU8Wjd510OhY
3TCf2vyQnQt9FX7uHgtMIVxuW10et3/wb2C/y11z/eyjzQSTSChKCfIgtCCCRfiZx2nP9Bw6lIrO
MvxOP9Gnwg7e3Gd99uTmymEGpU9zhzGwohpsg24y4J7dUD2Z5pSV8g777wjapNSxJA69Akfs9BYZ
RPq91y14il6vAYs4vcA+2aVZHNuW1eZB0CNSN+Q7UWrkXVJVA/1MSfpLOOjkCX9kVSQP08dIBiaI
olynIKJQW8sHjOq+bPrMTZb1XYwWZnRu9fq4dk3bAhMc3908Z3SuwLkhTICWg15TPjCOzUE5eYRW
I2caCBzMvi/HxycPQi71MveF9RB9x+TqnFJ+c9FjcBEqZyVdFgsf3BKmrXrKO5fX09/16nSO+3jH
zLHzvQAejWKXqTAxrFSK6LWqOWwYe8wxSC24K64Z21lIzI5waGf1j0KK+g0yh5ccXALsizQzk93B
VgZv+7pRKJVYye/pXYZcOsvqLC7+rX0MnCLtJ8yUZIJSgouKAA9RXbsLCEornNrOLtXW/f9o7atV
ZWnOzp2d4YSMNwRTRjtsii7PNh9zTXkyLjlgMm19lfJUw310S1e1L/H83BWd+TR/0sBCwWKuSjfB
MM0gpxyW+z0tFAFBE8D/hlvLs/4kSHYHpGwKTSUfnrh5Aa/t9GvnRKT2T0BCj0CDEycPmr6kggAU
hwUKnM3z1fhGjJX9kT8djotDIvlNto8iY4diHyf3XA5dbRHeeD0R9YybgKJu1qDfDRpjCyyyoFqv
3mazgUcCI7iuL5rBna4Uv7ivA47zSrhyDLIN++AbXhaBphQ9URL3an4W/eB8Db+Ck79ABMguYdHI
1+MNl0UheQuk+29hJoIEAk0BuO7EixaJgoH76ZxjVm5CsLmWLwxEiIfA0VuWBNmhtez1/HwcUeqE
+6zLs+3BENmcKpi/81gg6Kt9Gp6Jpl/OfPHslZuiMoQc7AcXsJ5ONfOmtGlXk6bZwjbuWBO/lZ5e
qTwlz0ZskZMmJzOMquXx92ElyIDF9dSJWkJcT+zGnZO/vjjdnONWWMs9+zXy/g1mm3oIg3csEdNO
E1qiAOH5h7Y59iyQr1KKWscf+YOBErDNddccL9lXiJ0qjjQOcoBQA5Ph8YhnUpVw37XTedDBt/f4
GicZPbfPBgz6Zphyb2IKh3CjGrqHtVGKaMrB13N7oRkM5MkTOl74Dil1trdr6wvSmJCDmz0Gxtzc
OV7X/Dgu3uNkC5rkyDw8FCro9wDmnlxXYhgGgJJGe7mD9aRaxLmL634rgFNhs6rOoGYpVeqvqyZX
QogV5l0pNHUQ0WmKa85DpK71zoKNeEh3lveXRE8spJt4b0GbCSzOsTjkBJEqdCEDuo6hgJ0XHhFA
AnOovytH8bQZKSQsQdJTzcOfAPjQ6L3SLO3XDxjfEdv1GO8GmTZI8xr80PBwf4pvJ6HpdZie+fOC
jH42Orzg3e/mesob8OwO7teYQVmmKrGduSHXkgB+5NvxNitOYx94fG2FVnOOE0SD1OiVPG07cndc
T18t59xPbAfZMn6oZ7Vw/VFIAZnKL9HZtPorRsQVxQG37XHqqdn9ktuYPI8JvL30uEimgd3TCUTv
4LUdhzCZB+CzI+5wLqTL8bXPLSDBqwFYN1yrAFqaeirMN164UeN7kS6t+YThvhID7Vg+RjHKAgXZ
9fAdD9UuieoPSN36bMaQTwEvoXbVfKKOT+pkhlYzv4XJgIhZYuXroEL3+VV6bHeRN5uaG5/Q3QpU
vXLtHooAJH9/y8+fX37fehYMgN39fZ/eUsuum0UoUre3NhUtX/0940joT+ymQuo+qdZwCZUcdEhx
IvbzGuNFFO1BOMapyeh4dXebcsvAHkqzCbYjWZa+VjWJoRsP6MPkx9XvdIAxZoUTNv/+SSAH3Io2
DknFdM/sRQ1JLkjXdGxpcWmAnUWsxFZNyL2Pp7DZs1PpOpTEdnNkiy+EVsTVYhjsAjtUQ6mVMXlf
GOCHSkpeE1Iz/k/iTkn6BVEQhZVn35Ju1bJ51/UIDPC/LZUzgiDbNT7pJ+EIKxJNrICk4bMN7LVI
Dm6ReKVHgXnJeZUlIkF6fo8ZFgxK1ePHSfOdbCp0DqeCyQgadvq7+qOxpJ/1g3fdi1Dd4xs4G6eJ
x4qmll5X3URePOMkFsGuqbu18AxR+81gHtznmicOeR0qFDy7uMns2W30EB6m/A90XiK/8aSuQYcz
zx1PbgMePeKhM9iOAD111hzRnjhTueRI1Vs9ygyIs4OlfT48zT+ClWW57kERR51nqo4MgjnzZWtC
SXq0CeDyECLywG6FlYr+AmkhNocUWtLypCO7bzOQnfa9u5MaOoc43SabG33KyWRn97E+653lvhgv
2Q05YJpX+hrXGKsQMqM+yHxdtadaJf1IYkmu+8YJeVHn3j2OG0n/RTzzLjP9EnUljrnwZ7tIOaXt
lK8OaV2ERtM8sc9EcU4a4D/v5jHjg3DBb6BCaM9Kj9a0fhnFPf3xXDXoYIAxmmZsVYWiBMcOihXF
8//uc5YLEqJ9/Zk6ppKdGsUs/EIzF/QnG2yu8Ri1+PbB4PlV9+S4LcFGzwqYwWMIZV+vTUZXNnoj
l4PKkrqvX619HQt8u0iLZZcXHoMFfXF8ZxRajHV5H82gxUXnCHCEUb48mUqwqV8/dpRorZnZUlcu
5JIWrLMLcJbJMcaEDMFduRs8pf6R86ZqHiY12ZsQqbY3WVDmAjHDipqVXXDrV2Cs9TtoGAattsyw
+arViqcsVf86ayXXUNVhdsdvjAj4bBR+06ZtFL+TaZPwj+CebHCAgzK6Hp9Olcbl9BJS09DzWBKI
3Z1qOMZVTqFNOsNkAI+sDby+pJoXEJ90L0c8DmjPRnGRu0ME0Ft/g7b1aZmyPdXhY9FGADeH8VgA
91s3yuhnRMbaf7em1p/ZjP8bhy2jul0Rk7VODOSLeQMm4Eq1AfBKtkoNBUmY6HV5nieHY62QsXXN
ShbDEbq3sHa+/P4YjrG/ShKEtkUQX+Oifq/RZKZrhvzy+VRYacnmxIyRf+N3Q0LjcrMX1tww8SxF
4hp9QTE+edUSbQET1z4MLwwYDmhTkx8QaSSV2XDzfRs+5mc8W9BNo61fYLJHcbuvitXIXw5jZRCI
DaO9huxRZUel7bLRZZgW8AyLRC+ckrFaTYz96sM/3zSGzpnzpX43NapZD+9SiMKRR0Jc6+lK9mqA
z5jFzOBm5l2KWisaY9oAgQc1imJ6KXFH5vTmZ4dmt2SprxyeKSKEno89cUu8VbZhmFLP08lf4DdI
5M34bGCsEMoltkkvYJquwf3k9bj0bXMG9RfcgiqFS7Wbe1CYsx4r19C8qFd1Vicg8f4noIoU+jIm
bUNY1OKqRyQS0oOI+IlBvRbZ1/V2JrVbpn7qb6wB0viPigAsKYX8WKyecfLyRaeUDW9YtPtRQ9it
ApttNZodoku9xHF6bDQP7rrfhWVLMUfU5WgSQFVH45sdXvJaGVvMsFnl+A4E2HTJ3XIBrsR9spOM
TgPEkAp8CLC/hRyeeVtYdTMpxGxrbm1sgzGxHj3h5V5mfj+lYt7ALI6SpjLfJAp4boO5jlcxCwsn
Ax/qsGEBk90K6n3mIbNRfv0CSbGlcTZTJd2VlojZfHoeiZbX5Owmr7nn92dtVfF9p5nML+oUofYl
tm6CiR5hCB4mnB1DIx133kGCGY6x2SsFbtOivK1S/6o66ogBcfgcwyL7sXDbEKCn7Z+7+74tCq5Q
YrfMIxLIZIlpzdJbIopDNlijUKw1oIoWCBxqz04EpNpSBeoB29eam0AB1Dpl4YZpE6eWSIomdGV5
+Zg5UMnyNg+iLIjQfOFmTH9/eovNFUM6BUn7NR/pUFWdYB3I2Y7D5+N2k7UCyCxYMvjfsuWIIdnM
pRgjXui2PJd2Bi6XNOZbi6kdxUt6DzZlubquc1DDV6hcf4pJ+/7mmvvRwMqN3NgpuS2ffXUFecP+
GMW9NM6DNlTfqk8LhxrWxg6HReo719A0ltGMS/kSFQmzKUlwVSNkaPkCC4miv4gL9ie57r+mMNCP
lmC6CL+0JCK+0xN4VI0+S0XcBuK/fWz0hkXg/EY23lk3LXgRIep4teQz0q00v7nI32A685Wxlev7
ZZJp9E/xciNtgCWg07zx/smYlWnrlSgDGCc95x8CIeGm5lKnuSp2IaSBwI0SecXndagjyiSu9IlT
I3Q1FdLbg2Wnc7NJS/SBS7gvnOEdSMa92dsEUf2Oi6hQ475z0vAG+Ep/M5b71lelDUpaHU2q8MqZ
F1slLn/SnyLTjVvSAvv7CNH/Vi1unrxBfksl9DBQUHKHMHn6k2Tck6jaQZIFT+xMw/BXv3Vy+mAK
sSjsd5vH7ddSpTJIBeOrSkN+XyNSkwrgOMAkZtSCqPh0wBlxwDPAzFYCLS1VL9sn26q9ibve3dwu
zYwbtaw4esW0C8xskiDtgeIFE2QhR+Yu9gJeHRCiWcfShdWuGxxVlW278cMeJXFv3DydN4WmvcTo
QkbFKmi7MUeBh3EmJvlqFel8nJbRLNBcY3GJUlDcfbuPXWBuPA6NnBgjzyJ64atngeLw/6G/Erx2
m+uhawF6OIMrzjr1HUnHOoDbLAwca3XbFyIe+o99EmwJt4qcxcILxMfxt9YrHK9QyvK9csHkxzNL
QWbs7p3a2OhQq83iNBevgedmsXqUv8g55o4uTbYSe4usQzZWNRk4mYdrhCdIt0fmgWKv3e2gdHl2
KwgaxC2rgym+rTsx5lQ+SxKne3IDmpLrFxrJFYhhG0DZvmTlq3kI8yETOC4OMpU5ep2wkXJBYSrt
musB2cmSgbw4x1dZ/sfaM4CZS8pF5PvjW5It/Ato2pvMl9CHJYVde9lA1EGFIIiSdWXm+fRhZMw1
WxHkgPlSbcdj+XSrn54STG51XvZYv69//DOs2QW/c2lsBz73hgq1hUP9m6WsmVZMOIi1rTWNBIXP
MX994NGAupz+2UH8WN8/p7tSzlapcHdc42fH5ST0j+D22Zrxs0eRGe5SHQY7oV1T/beI0CbG+L9D
tFXi2hzThAsFLxazmNpVENy1iunVPDkee2XWY4PjaMR1tjVC8Sa0ldLtDoNm484Ghg3d5OtUxeKa
C8stabmT3PYBdf61+oTS3aqF3CYmnQJrTm12sR91YdwqlGrYPGfdflHBXfxFA6vceJhKwGKyree3
I0D1sB25EqFhIHRBK4piksqFwyeb9jVTWlZYpVHzmhZnUsWxl4ufwxumnECS9jW68EEYq0RerhJD
xqDDXbZgs1AWUtCnQDUpgVXy3Xtb8wBXswwpXwLwa3TwVNBBTvFqX8FwyPA9vxw2dCC2GbF/Htrm
4UE47rakqsWOAt5Da5o+wbfz074NDsDBqDhLUA9se+29I6Y9dwX2IIC7GhgP3kSn8I7SI7d0A2gZ
dijIQP3GzEvpjZOcsxyMUppqM5zMK3ZL++jG9qGnMz5txirK6KbQD3hIhuNlJjS+itG84L7KQbjO
GOcjqeVrtnUBY3Ngqmnmf342CknrNgfVS7jmvyMFPw54+HhsrkH8VbSShhXM+5p81dZqNwIj6scD
vXsCXd7D2Hievekspc1YBvQauV7LBtJf+C6Ytl1ur7SaBvzQ2v8boto2IQnbO+k7aDw8HCmqcTwV
g6zLbmFGCHpNc1l+tKY5bHXuKe0QcWVqLCQ5gBWh4DBx6ZGL8/zIYUZhNOQsDPRf4vyMGZxnKup1
/jtvKUxGRaH+1oIjjtjpndx+qg/Y3EtU1njMXYmk4LvB4PJjb21WxEyu633fXTYNJUc+0rMRMlfn
gJnuADU9IXQtjR71hKSB1oGP8e6O+D9T5QFBCdLahnSppvoVCK38hOG8K0dHEAyqOayJSV5SfVd5
9XWQdfrFQrxXn0bICAhw3xjKVCTWVtNfABhJ2b837AIl87AGgBALfuQ5M6NR8ZGu/TvwYFsAyJLC
wOunPkWmi3fd+visAffxik92cRlWWRmKLwXVzOBzxnn72XrT9RAmW26yjPOrpdB57b/+MlLoamgx
HfHFO69n7xWu+SI1NHwRkiDmH9EXS30cznXnM5s6KFlkK+PN+4BYMitsblG0IAIeNnsWON+4sbZ3
dUZKOeW2d7yV152mqbCPEhX2KKNczXJt4ga8ygUpcaONNJT/7vfUHrZh2zXMVnBV2huzoq4ZFUqL
JbIq5vYiiBKp4V4RjUr1RwhA8U1pJMoe+v2QmhptvW9ugqYA7ACpnSb5yBY/caaSztp94QlhFR2T
SZ+D7QmMTA7B/VUEY6tklGagPxPDrdokk7HFRu3FsOK4PX9xcL8QaRgbYgPIlkmrapMhtiMNsqak
lA11X1f7EY4bSvDkKet2xvidYvfpTiYQHjPtV+M7Y/CCGWlUpgdK6E+hXF5r3nS7sRSV0/PdV1xL
VHd3WIghGQm+FEIY9ihb5mZZNmiCcijXx/LU/Cfyk4i0xZch+/9+YBfJOc9edRQBVicXe3stYn46
efmAK1lCkY/NKxbD2SgeM91XHXZl5CSdu+jz1E+UNQGnl41EsvGq9iPayVgFDsxUSlLWJk+l8OxK
bJMIt9bGOC64sKcl4pnVgX67PfwrCPnbzkVtxtdmXpCpz5ivTV8FZfH08Y7P3HaKQJ3qXTkguJFr
TFlE7v+bzHSeTDZiblAxu609bDdoLPz91uaiaZLf4wb1DuFaDyHsxCXNv8dk2eC3W/RYt/IlCK5u
1lWTxgf9q80Tvb9/PgAjwe/gj5UzaBPrLM21C3L99pB+SNzAv5PXCfFCn5LfEsOpmd9/96WDo15v
HgIzqGuPg3xqVBb4iVL5b8XzvXKf7FLgFP/UpOtVN00mMFRMIQl/Kz/gEeRSVGtiqRJTaDwd47dR
yfq51eLIsD95MZErVWx2JCh8SE8TfgwVhWgBPFv7focxElgiIKRCB5KyWO9IDAFBEQeGM0VVv7/E
VuhVNz78s4f838/O7CDPkFL3xN+Bm6aIGXzIKcZeN1Sr1n9ZxO4tUceoxSfis7Xth0W7QNy1W+4y
zIpaAn0owR5Sy6RxVBtg+jcnb4E9DI5gaOvXfcmdy15EAmL8isn5NjFTmEvIsmmzmTkroopVM8JG
RqRtBomQzUOeVNbCVLl2XF3RsxIXUKjde987dZfXDB78Iz1kPq+4W2BCd6kxVYpMVCKm7NlyhjTa
vRxH7c9ub1GWgDBoB8kLRxchypLGEb/v2k4eQfUKpuHS+i8ueQ8A1Lk376pCwIPLDyGkmSlFAkOZ
7E+XfrELmKeRPcgM40QhjWwiA9Y3tb9BqnTe4jVPbJH4jKCVAtTWkHCUipRV2Am/v0gNU0ek0Zbr
T63OyBSWpZp9SRVwrb6hOj4i3UjuZC4ToceCZxSm5tyP/efmOkv/yWo0zrUUEULl/y0vHvHrYtOR
TYl89ta0ZCENNWUtpKuCtGISyJ+esF8bOYnCxRwiBO2ic4Ivw5oeCf3vnDnR1OWHKLZ5stCfhtMd
p8oZIrTUuE/hM0W3c8+S7Qx+BfGlS2387C0oqenwZRMB43bOGwpZWiVatLIVSpA2fMnOvGO9B8dd
klFirOyEsawg9FeD5sGNOjEZfObdMcjfULTOliEivsnd5DeAybntkuHeGaGU7QQ22idvQJV865qT
TOq07/hkGdMWwaQehQ4sEqb05tIt2UJfdxbMVr09ZPOLjrV82xiIgLIBjCE5UsIZMIZyrxdSca/J
qGM8+wcRNGHk88aetvdiD+m1UgAOze8h74WJivDvJJNwk0ZZfmiChYOS4MSwfwG8LqT+0WvuWkET
7BuELx48RW0tpBmhGvH7oQ4aJiqYm093wFS8zWZJcSlzuHiwC24GEAsYMSaZX1F3LhKWA/VXsQsT
QJqK4qI3jDQvLbMro+SNESFa5sNxvghHCoFDLqpXYULtt7N68mwaic/sQsAM/V6r4eLFLT5w+pK3
cM2EnTZKyWEQy8m4AOAqdNfrYw7DbO6jd/lTuORJkYwzGxxSTWVPjzXQBjB1ZBxdnio+1vx7mve/
K3wvi1T2dI4di5IiPej/2IfE5Cd4d6CZV7iDUQBWJMTgZOG3913Pi7KwH2er/klorAUS+fKZrzP8
J3C2M5lFe5KNHfh+BUaXJwyw4cSCV3i9FuhzNhCYqyMjuhqpVWPDIECksNWozKCvB1aIqlyvxDQx
T2TWqrtGpnYsAMCsIfwGpMGbyzClPN0JifB8qAtnWHxiIo+rrDdxmOYmSOrXgj21xKYHvrP5Asku
QRKqW1z5Lh2q+VAt+4ZY4dLV36tDsN5YbLylbcm2w4m/kVazUrgygleD1SyIilbg0YuybexXdzot
Cz5wd+AKvR4W4zusYmAgO28LoMLmQu09bdlRpYjpOi63+8Otq1E6YHncfnf47nkMHDXzWraEwcGA
fLZARBHFurUsX9jXGpW4tx9LdXPnE5LO3dTxAa+dGCEtU/+Rk34t3cldM4x870FQFPbGgyN3R57d
X7mykA5Ck9dp2utUEets/S1CXw2ROBS6NkqsLG7eoOdcMChNi44tPMVeDuBUrS67zhW7sGp4AjJW
awOg4LuRdrL0dBduCx2JorQ3fGjFRHGmpkrma37lsPPLrX+ZN/iGn/AuCs/sSCwjGnctoPzvnND8
AqJPBvt2NYVAjBoU2ABWgzqq9YzLBWhAZpc8cc1iT3q3F2fMJ2fVfJ3DtfxCMQTyRbqKGzTzU+N3
nq9Zrq/ut+gM19Vm8q1G84ZL+Yv4Gr1/rsnnoyrE7x3xW6ANbuyMEsND0kiPfm8p7u51RwvgAToQ
H8v2McrwnVXQFe/e//3Tly48gcT0lcaN8wXF59ULXuhXr935iEIjCA6ZDwbipuRaivkwfnVvNLJp
HevWFXux/f4ZBip0ZE6/UeRhF3fJzuUiEVzLAND3PMSO3CqJoxe7STVXu/eyTm4CJQNXTKMVz5yE
WT2ZvFPmDVsaENwr7hUUv2l7u/kHt3RVVOEiyl5lS9viCcDxAuh0DQoEeKGxZhkJ5+CU4P5bRKgl
aLnSMd0P3rdT8S/kI2Nu1wxmRmK4bBgNqnWHQGzzAKAisG8+wsZJ+q97q6WJRyaxOCAkVnU1kJWI
h9PJGfoPJRozTrOIOPUNg6FsPA4RZeA4/g8lg85qwB61zOU/M4vgFggOJuHQipF6o2CqmDgNs/DB
cPh0rbuHLSdA8RNudwa8+xZ8u5uRN6vSGxfDdpxh7RL8maOfNKwUnzcCyMHdEU4KWRGFpAbr07B0
q6aTaO9OSSolgTbMwr3bBUfATjeBCbacuVuisxbCcPPL7EBM3Sk0eHfxgBROHvBJlQuSg9AUw5Hg
P5DKG8Tpkfy+EbbBxZCCutZpaS58jtspnba8Y3QjjcXH22kmglwPF58i1ZEbIu8zgFJOoHgzELHV
FNaHSIuA6264e/gdlJhZ5ew+qvaqxCkCyoMS2uKVuEfCZZDSHNSi1qJY/tQu7Ggb0JbwPvFKcwDA
d/cZu5i2kBPZVhgsCCa9bc0UGuUAmgUYGR95v7L1Le5K0Ohs2KYdRUh3/pSBx8dZCy2Q1YbiVbF7
M6Ao3LZB6Xjls9yrAf/ls71j/X1bdoH6qYFaM7r+6PzcIOQ2DOAg20pBSRqhmC+GqtM6Sy4Q9vir
4mzEY5IT0g/JjWz6UTCpbeGFkjHYrbCYqf9CPsEsAmJM9DPHNgbODfueNHuZnunEdCQrdSFuw3Jp
RL7u1VhVj5GUIiqe3BDftVS7jRXeKbCT+yUFUzZtUyVzE0SPL0dJIvor+t2QIUY9M2ewgFkIQI9S
4tLcOKmMat3CxfZfjeEhbEKDCeBJm762VkiXBKbtJmJBvQHF63DGAQG0mxEouZX7xfGLufPFsdp+
MYGwijQUvgWbot/dyFxu3kfOj5Pjn17/S2NQf55OwkM+61j/LCrSig0Rx4PfJaeB6AB+oGDAkEwO
FagDVVA6VHMqNu/XPUezDZl96k4/gopwk3CJOgNamDEHqx8kI72ZEgWPq3cK+KFulEZQcRBLo44x
E5McK1wQ38ZR19nKhQ1lwZR8/b9kAMDkwauau9Ve22pZowxULSc78fcz4jPkVS8cmW7+FIjhtG9P
WGh8snraQH+apbInOxcQkRDTzzCLRTQ2VG9n7LaVYY574PEcbKBAaH1xoEGTGWG/gDZzkETQjt2E
oS2H6wpbOtKJMvhrBAicMXmcvTB/19AT3LHRheuc2oi/YPBDO3TQTwbBsnBYp5Ktne4+P6DkjNpv
QqjUVc2vZBLnj6/ybNYLCTg3E1tKqyL3mLInXHGI4vutbNvPBhqeWF0KM/IFt3WXDOuXUz+rBPfx
bozTStGXR8nl0MfNltfi9bRisRka4A0gCIVdQ3OFjTEOYS/aAr4I7bqe4Ng/YpDbWnA0aFq73q9f
WTrEJ5nXQYnpqHk9HgiZmloDffloCN+7LnRcoZP7782BbnIb4Q/Apa+mXYt4WBbfmRMrLQfmA6bx
KnVfdEFtBNeJ/OAAXOBONR5KFg6/ukoWcqcT5Itu6ew+2nXPaLuyd3b5GT/2hvJJmU1t9tzY9Y64
Tx2eHxB3xS7PW4OS4JsGI6j++csysUZECe1Ctl/17LC4U3ko7toB916oR3oMCiE4uPccoMbL2R+K
ewXhJBBW9JiEafqx7uLJJJMi47VRDNEB89k+dI+Wripr+KRhk1Eg6XsIwm40XbLHOI8QXS70G2ST
FgrvOaWSMGOaiaauYLA2MrnZTOhnQTc8bgYFflZUf09lnlvujpreK8s9I2STdRnvpNyAn1FYmwUF
7ubOIePAXlpcxdirLHDcElROd7DJwWHjL5gVfjnuimFnuBfNBsPliEWKEMqEE6BvX3kEtOdHb0ms
B9UwAYr7cSMuBKQGzIs1my3sfvTINFFG2q6fKxFuGx2OVFMCnj2Z3glfJqJAJc7E4WGfXx/EI9Dj
To5w5CJZcw6K881h/68O82XLyAtUkXYWndg0/SZ68jdLP3bsaFoqzyPva0KUNcFLnHAaUu9y13A6
UJkrLwWXKPUd3coz9qQ9H+0o6m8m2cNUW99QFhkRMlGxjyxfvuhpSfZmLZeBwxa7U2alx73sBE8Z
i0QRvq/W6oVM6E6UNFq2yJ6T9N6tAZYBkDDtCUBFaR6VRRyxmBzg67Jp5ILT6N6LkshC4ZoqadJC
pU4PiytZktF6VUyKqps6msalGC0Us4WF7sYr8RUQuoxZHp07hTbQuAiRuagrKF5kQFalqLzk0rX1
SOSABKnxKrPm1FiPb3EzSmOx59PQOgAAnlggSS54woEsT/o20gOTn1gvUGNJtAteymTTJ4NEJ0Cb
Miif913/AaIMUnlurmVtq+uIXgrEYdfyV4SgsHXN2uoAlE5O2D99kQ7NmDoS40IvlcjZa5MKUExm
dYulyR+c1VpD1hNd990Nd87ExjAYeLW9WW3mfnPzVnv/iz1OPNlDhkoT+QO0ZMiwb84iwZrT2NQH
sfvYSUvd3GanxU7++kbO7i4s/nTwvtGSl1SAb7cqz/3YrSKpGfldOSwruklcZ49YP3WwZVo0sf5Z
UrQ2Sc6ZNwSqjxMnZFp5MXlG7ZVYVpxtH1UOVlTY6vdUBLPvYEDrjv8yH1uESxO/qDaHCXS3cAbZ
AE5QtrYt/N32Hcr4EWoJ0hmh3nTBkMjidpWI32AYWRMDSbAOQcmfM+yaK1Nq/1cuSV2TqnoGfMPP
DHUxxqgOhPLEauV1LnrgUFTu/lSsMLIrWNDyGKh8giK0BVPT4YrdljnZAW+QuVGtzUgxfY0FQLHH
bROErO0WnT71xb4bm9GKTyctA406DRqnLkwAfEgW8I29n3J/PFIB8DQyW3DnFF8GE491Q3KBc3Qw
R5VjwrPDpeng37csNEQ2OBeXm8IA0z2GGcZLux4LSD6nRVaFbrdl1RJvZBiT7OwNi5duiUv+kHEe
LHcl2JaGPBF0rfBhMYAjY3i+HYJQAdPnl+Zlt4Kb9zHsaUvQSFycIaw/oLxvvXHdoYC8F8hPgfON
Q6pnd0XXa9T53MmwjZQuiuHJW587c5PE5txslYwSsw6yIA9U+TR8+cjNwc27ZN2XJ3V6AITexWLt
sbGM3kI3Xxiwp0yTGtD2SkUlCIIqpl1jF/ndZ6tL7rrIVVFYBbxxLWgxYJgBUiY9Vx1Urj9LXbK/
MidmR2F/W6h8TZtqXExDItRrkfDVFkkNF78Tif7aAvmpmqCjBFqk5LL4hqVzFp54czaMPxk7WD9r
MjRlhVcHcCjavMWSCRc1EkLDuS8cyGkIP2ItQRAB3Y/Phe/eFRfVEsksefiCcYfobxyt4OYwwSlO
Dy+DYp2vTVhY+QK8UCpH4sHxTd/EQXOPARZFhy/xLWPochyuKV8w0Ygxb/n3xaCjV9x1AffM9rJZ
6dq3HRgEzRrWWueR4nFxpHDc4c0yEV4UXLXw3kd5zyzVUeqI6bDna7yz6/G0NA+yaBrdJ5yA2wgb
R+Z/bWudLMAGbbeMfGY0IPBFak5Nq6u9KztuXoGhH1kUk0hVY3gDPi33292KvJQlvmddDf/uIKKP
bQA8iexU+BwOesX+/+pqrlMM1UySdBkwjDDr2ytrTif0r8Krhm3tgVOEXhIkeFxP+WALgaY/zlvY
QfHQcFFAwAdSpj2xHik1JPLroD0qQz7+Wogqh0jHr8WFv/r/baMfYBh3PkY+MAsmgcobP6SeYVMV
X4mKRdxDPKC2U9egWQvVOb3mdCWZTuR86jurryHG3+EdKEX8/JGSnZTfEuWBpHgEXv36G++Q0maZ
3j+/HDe+QchzoQrilosuZynLi/EFskAlNYoeuUPr54Ecs051nhDOvp3X9PLMYEGwXcyoWmBG9tyP
SEL++r4/6dt47ZMim1tjbqY0nOjWJ296qB/F9zO9rK0js7TyUwb8T6pgoBDniipUhJRvceqp9wDu
Fpxuhyjq1tbvjoj9tjoI6H44qXSiX02VWMfRPMX5gjc3GvM0LpThuc5e1LP77+4SMxtVNGBls+lb
f3cYsHsJlghD5Z2SlAZzD2bdTGWbYOukHsK80acC8oz+mgN/eOIt9Decj9mbFgFjAVUvmJKLMduI
qbx+olI+itGr/MEJCI+W6t+OJklr/t4uF3iJFmqsxconMqNBZn56Kdtz42kEPxqnoA30EWacKbLV
5X17hYrD+BYT2c2t3I+93ZHMfQCe0Nmd/D+vCT1z2ntBCICYtT/brBqonNfY5gru/MuytSg1sPp/
ugwYXc3xc8jp6p3AJrdSDf/rH6OZD7YoylOum0aONUQ92vcPm54yhPpZtc2HwrAPLHRXDNfSb4dS
PWVmocjEktaZ+4B+7MVjjvoExWm3TqMkFXTpx4JnGPXRYZgyT5JLNj2NKWVWPZ6JJdi83KpkrBxm
TBCAIQtJZpG49pE2nZuGnirY9mqtXkoT5OW5E5U5aJO/YnmhJTYuw1bTeaB1R2XV5eTaFqjFf7eM
4hNcOIultq8lI0612KR5EpDT+jyN8pCSu8Oh/7DUw2mWAfiAjcJWO/9zTuEE4FDD5zQIQlqmYCwa
8wg8zOVRieTZj+dP9PvPtqsNedWOq6JrpHYBryyQ032ZYr/ipvxD2PKoJNcufbM/HjyKbC8dFugN
Ra+Lag6cYRp9cXIug/eYB1H1h7dT3ggCcTNCPpER3FpeWoh3q4eEaAiycgWTqJvchlv+BRh84uId
0AmYJKLqmif8HvgHMFHNl9sjXA/Gn2BBUeGUEzvG9XUlPYG+dQuUq1OygZQ9OoGoTc4ADcpSNoxx
kAUxCMxT4zHcbKEM8dOZxpHJXzTo3K++ZVNtmmBmuXtRNXDR1XbD+XZqkbSisPc2MLGKLrQESjiX
xSA28q3CmXDRyq+rqUGagFC8DPV6IujSWEM6U0YQFofSvL2NovTJ951YsvkXp6GRA3Cf7MgEBb1+
gE2pC3AUJFbHjokk2e6+npFt1m1BHNzQ3c0Wwqbdr/0yhAkO4SPQt2Kfx1IgDK6nI0W/BUVKQJcy
pvXWbzECym8DY6QWJ+qCG6tQcF024yFBjb5A3+z2XGgMoWwhnElArTl7Rtm7VC5YTphZ7tkVoVVo
iPSfUTPzYcOgQudfUGGqn9BCsdkRlaIGm6FqXwJzmnycXabYX5u/b4ZPog8A1Df0GGLUo64HI0hg
yybCNFAK6IigSgcx1BeD1/1ZYO33/A86l9oPp6PPqtXAMNbPS+6bOhg+hAKy2cYb6O8nPDneljzZ
dLplJFwrL0KDw/ojd1QpmmdRZLhAcQRlETRVcfinhwQcqeqDkRqLiqIjMVfq3Yk9/Y63Y+6la/7i
093KAm1RLQNnlJusucOyKI+tP9Rfot61c/cEHoz+VeW+68fZV8k4qospyYpivUbqolB/EaYN6vky
L1Vj69CZ9qsASxVZJjrKO/U3OQoDRz+rPb5I5rmi0l38gTVRk02TFVe89WW0uZv0W8huAo+ekyGh
jUT7vYI0+Wrgn+n9IbA33woOoUrD04B2xnFv/mUR/uS/lh6Vig96MwGRPhJMcfppnQ/k7GTU3zH/
7JJ392jCZjwrlGNe0n90WdoP30KubzwS9YbXGuDMm6328ph8YbY5IrpwJRBXn4bYmpZHzf2sbFhR
oLk3pnR9vrrAbfoyEOj+74dChUhiTiEA04JSV6wK4T953pYtNN9x7Y9Vq1tvtqBBqb0zdlwBGikV
E/LVKP4rvhsY/BwczI5sq2lPlO5SLK5G/ePdherTeiDJ3A8h94++VROd84z25XT8YGAAgyzLw359
nTw7LR3aZbZRMhVsJ9fXIl+QAaarw9MLoRxR9jmrpy0UWAXOouWjxpSyNHAajBwoVqcpvUAazQde
wR17xoZk4Lih1kshMmWPBgSLp7FCqPjhbgYhPhzYrkuQ3Gn2xWZmpuKZj/zxnFaADzlWzAFaaztE
gWoBn5jA+4P7qUcyoa/1u04kY1kDL2WbMkgmvG9+2alID95J7aXRP7AiqQ0ruDHbIY1L5gpQkXpS
CdJqfRGDPJy8bgVIz9YcHbS6AkAkqfdMUmcH177BEOt4xc8U24b7J1JXq1FSf0C3xNMKWmDYlaya
/bW7Eu07jeVAJPZd60W9MsDirZz6rKqDQnHpMmOUeBK+g3rXpjdGaRf+uNwjklkR89wp4OLN/Eaf
tC4dX+sG2TQJRNTwbn90JmNxRMjmCRDZZ6S5LhZZBD2zmZjEjHHYR2n6ZlPDHBGRhZOPIM/nwpHI
VbbFyaLCIHmaxtTFt+T8366258nV27mUCGSzBq2CRI77AJsQdZrLEpdN/T26llyP2+NBbShQnoo9
YMHhpUEH02qkMaCpb7NRBujfCE6N7+qLpT/KATKb/aAtbjLqLufCPtolewR91xZ6h1ir10OB3rq3
2HEJAiUBUDge46tbUmpAYNYx6ke7GQnt0Y8WAZ8zD109HBKihq4Tzpowk8ejhvFcpA7/3tJPiUbq
B130ixPSxTvxKY107zyIOko/t3M93OnC4GsAseMT/ULvCAKVGOvoYVjE1Tlz3li4qIwgSuMVrS6t
V3TxGWmNQEDVQq6sGRhU4Jo3Q62k7N/wRBO0yKiRfiN/0exL7Dua6JInkbsaTmQxLlopaywDk4gQ
nJFIrNPxHjnhXBaMWdfdmR6ho+ocAtvkEHdIScqfqJ2g+IsXqOakeV79DnNiwU7u39/Y85RZNyg5
85I9u0MU/3/00yp6mndyxm4rSgM0wajU0nqxzhZFwi0eq0fuygKnTDJXSmX+1DbDo6hXJqcPXoKB
xUNRhpH8C77n+JZRob27+XJbqNlzcrReWGI5nYV4zNZwpj5LCiF48TlOFdMY/oUmGf127DfXIeH8
kK0IAlN3Ok9DGq/vZ/E/tS7LjdVZJ9t0UPltf1Mi8DSs7Wwuh7+kP0ZyFQmUcuEC9MrITZtimmKj
vbB5rKDTtqIguxHdFaL+j2MO9GAyYGDjkrXAYYVpDmNCW19XubNunOmsAVpLuFsPxtg0sLFagAgT
a8i9I2Fmc81Y/g5e0V6Jh365J4KDiOULajTkWrvdWq4fiJ1zimH6GPgDFjFTAby3PnhsOevaxp9Q
20dYBwlPv8Eh1Om7oPmtSKnX/E4rb8Ly6UmKmOx8Gj8LxUy6hq/C0iRR7Ll8LiWvRRHGKGt3+ZRh
2z4sdYWQ9SbzFRHp3pgdzpRECTHQoY5kyqwKSiNEMYMTShuD2wWdNmFZWUC/DgMzpypUUJO24oZv
/+NxnBJYshaxZm3kp23yWyUKICsquD8IgNGmuPvWwa1BfJ2/3j9O86NQp+GkYfBoE5xSUKyRTnqt
C1ZHwYll3SooaknQAKjaGK4SFq/42ZC+b1+l1oyo+Vf2lLk7npfggr7fisdUAt1gL5TuEbF+BfFl
Iec7nZke3jFMLMvhjeyBLU8YQKn+GCrRtvpMVguYmWdqmhBCNKyNZEcr+CWmlrKFg9r8Tnj3J2mD
W78rcCXfjvZ4kyP1xSPJGbb5valzizUfzjoLbxA5eHSvnR66UNES9Tu4U6bsgCV128mz25VUHgm1
SW3ZdGDG1pf1YKRwhUE4pOPWbDLQJ1o96fHJ5Zv2IjAmz+pGJ7+6XtfK0qVhff4JeVS2uFmHKER0
q0e81Y889MqhmWVpSSizZj72rYqtz3o+DYjCrPvFah6qn9crYNje52GmlHsf5TRtm5tuCdt82ZzK
IF5FnMHSfcdLbHp81oo/iysULRvrvwyjGZWlv8ZoRoTFDbBCdQn2FZVGFLLcl58UeI1+3VkzUfe8
1EaUwx3sFRFAAHPmwGPko0NSkjMnakTgO9HHvaxtFkuPoHPE+w0KP7PTJ+u5jWjlbp4etcGiEhUG
aL3M0A2fRLQJmZEyu4odQgj0vgoj3DIla8Ub/RRjpKF+Fkrr8axq9AK0DV3RCyt7h9qEM1yWiLxo
90RDMCaf4rRIroGWhNK0klSKYde/H9DuJzQbL3qdWdeLQcB5rSZ8GDBhSoOA8btbtzbmU/O2T62j
xaiKnG2ynOR+1kclhLQb4Qe0J+TbLluYO8KICG5ti1bPE+Xv+juztq7gpw0Hksn3GCTeXQwxd/bf
6kl+2ddB00tBWQBd2ol/dBlA1tR5pmZSecno4VRwazo1kElywkHJbFALvYPV5Td36ZdDpyjObvwz
2F5iR5O7nE1vfgl0Bdvz+a1h1k/V6JvhRimpp6ZHB6scED3skHYcCFbkso1Fh9uCy4hPAKP+Gcm5
xC/52luZtJffSWXdzYJbWIYaCY+5budiLb57fo1OkcX/ZnZtuyB5u1RB1dRP3R5pV6iH9ucLRqTY
2MGcyctL4A7Jm7v4NqesS7ATWVhrzlI0udmf6LN6mZCi0H7pPUmO6MxA2Z9K8iAat96ru0SYe6Xd
RxINQVIFMErNQVmI2MTZyaBJIZeTuvkf1ksHUDC1yonp3vV2ppMj6FaZrBZNRmeawf1yrriarn3c
KN8AjOLDAR9Di8XKFaeL6XLcrZPB19/1hlEO+6W1bRlYM8uVxhol90ARxcAUjpZ9qPoTHJVQLRf9
MewdCMt2D3C0PI/LzTij/VQcryjfA+TokcxKF2iYkwWtI30CNCL8Pj4kUIsfdN9D4+KvO5QDS5UF
bJ7ORYOIk4bpoE+t37mON2Zc+gEkmMhDnCXOLoM03v6gS6dL5SLiqI3mmXmubYXeTXUE3Mg88E9n
CZ8f1R/zZ+0cmu3xuvwd3nOgkmDhhIJxSgRHuxmIHEbDr7d87jUzIwtT6auSRSkJdmnsM+9xeYtv
BitspE3kwWUigEJ2R22hzdTtv3RWv4iKp7Dh0vaTDoblj3NP7D2dRJ5k2WY9Kl/dEoD7UgvwxJx+
dPRIouotru2X/1rh4zgEEgHTlEjZvBELg8pvMjWkOEYIX1/fqnEN3x2Aiels5r2nN2KfvzZAzBhW
KZzPi8HGj+eZ+WvK0hWumQilJKvlAsJF8+mXXqBIfTB+6cyoZQWQ0M16tao2GMIRwlX5UeAwMQGM
eYIDm245IoU3pUm0/eSEqLZ7UgYv0ls2hiG61aZN0Kl+dqLCSLCpCAS1rTRa+TOyWHeTukzxiDVv
vnXkCgv0E8TmbtvH00oLwTyF3frnnlhWN28FOn3eqwUiqs+wBmPOnzNBC8aMb7T6L1haICW3QQRs
80Kvg5Om4JX+B6AKt96DtYxrmjy0xAYAQMNoyp23jvv4lv5g+66/asUGUWPFGiVWvNhNDNue6HlZ
jkVStROjq+7OsyopAXXpxopF5g7Kxkwxh3KVIgNjXSZqpQyOOk5e8osKloEYRwzV1hWyUWt5DtD5
Nen9uaC7tpcVsSrl5V+wnH58UrOutpUQLJV6FjJPyYkHrXn02CACTgiahGpoiQ0tWWUSnN9JnMIk
aTOIELHqeDJM2DRJZII3JyyIgu+U/QkOYcJA8njTaYoSjMOA23+I/T15XhHslnt5wiPmwsa3ptOe
0Okxz69ZeaunaaJw2ILgGQSy1JZ1Jn6wOw9YGqt7368iGbJ/d4iXivvGcVfnB+W5SK0+7B/885xw
Pnokkc3EDf64sePpPnU7mMfpomWgVI5DNlFMB5/S9OV1MHyl8WWfv/7znGnW1UHTT2Kza/1aXmGV
bSlcl4FHSHqRic85MJQZToUoa4vMchfiYonY6QvyJEGFtPlJVnrkClHnLbs7GK+zzRUEvL0C8IFv
2ApxZ33KApRt9cF1rZi5sBQIfpi1ozQWP32GeQjfThHhQeAOfscZ9ci0zIghx/JhlX9qWlGukQjq
B+qyQLiR8fGV+MhT9WTWzYAJyR2ErhpRvtLdxH1JKW/jjV6iLs1iUN1p7nSXYkHg0aG8QVeDYu1R
xaLlXDKLeSiMvGT/MzURPH+Xk3CC+gKuqsrvPqiCFRobXXa7PPTNm2pl9aw0tyqNboHAQhJ4fkk0
rsyL/4U3HS6zOs5RGuDorKDfDbF3KZjp0GtNBcrFCp8SyCwWl5DUOyxAxwNhZqEkTes0lVXyBvva
ILqekBPCDYu37SAIsPrv8KUoi+ld+Scfr9+yOn4DFSINynqv7ck/dgZsNUelBqAR0pmh5LSElLTO
HflZsIzhjfUbjzvEYFv7EcJPQ1MWRVwddkTp10HXcc0kxstNlyAcRlNzGlg0R6sB4wAmMOz8eGRg
N04WcFjfowQXUy1tF3bfUZpZFygexuNQb2kjAc1LLvdaeY4BaF3gjKzO6a+dO81kt40R6Nx6o1yH
Lh9jBFoyn9+qEIOi28RNhhXtqE0G/J2RHLU4BH2uq8A5kUmfpR4G0MZj0OlsMWxFMrpQUlspZ9sG
z1HrNH8MP7GwzdXUkcsN2i9krEWcppUljvRCdMZ5wHD+FVPkjQS5PbvcxpbIAAx1VxfXus4fDUV/
dZww+91xY4e/cZ5dM6/P+41ZQXeg2MgHkm1v68uNs6fgElaQMybWirC0spkbTyPgE+cXTZoRn82h
UGmsAF6tHkg3GlkVH+XyvvT1k5/cTnp4O+ydwsh+VEvtPe6IqzkBw2LQvxOdPQ+JgCi4PimQbB0k
J/z9Rg6WB7QkziIpg3UmxgRt8fWl64RqMtpaQsv3RU5lz2Gl5L2GFycQJyPwE3gfrZ4caaYmKZHI
1liMVh75SQ0xVJfcuDc85DijMIxVR0HbjqswKUP0tZ3QGzJqbVgw3Ozjlp9u6B+pCTiDEnqcYikZ
wH+NKZJD/A45IOC/QaE5qywLDQ/IMqVGR4F7hEFos+wxK3K660+0VfiEJj+qdTJuud9AeB7A9FaY
Kct3HHvP1bRKXUCVy+GZGzXxKVF+PK1s6oX2Cz0mbUi6XHHLkTTQK54nY+SyzrKaYSPLiE425jQA
G1H06VPYxm/vIsB66B+lOLk7XzlMqMw1FloY0fvyfqgQ00eVcsGOfXNhO+feoFLwryXR2BGNocZn
dLSpsow9OOrEWj4UvENQGWTOlW2TarcZTqZ6+FWY8/99f3Z6MacEOzItSE/Dx9aJuIaJXIOBCl6t
Z2JPHdBsN+gjBHXBzGAg0XhZeYi6W6b1yGz2Ck+juihcMKiNFbBDc4KspVxs5NQF/vXwckOQanzE
UuonWd/Xy5rbRKTDoQ+3QVmhjrOWBAJ6WTzLkYkhMj7DpIOXtkNMUnN3Irw9KooPzBnYhRYWvd65
WQHF4GM4/on7t0dmjVhwB812GFgI026ak1QTnI/dOeIdcAJrX8nHK4QGoGryRESdnkB2OLaB8rAE
sV1ySgSIB2E0rXANQgVqZ5j4eJ49Fq0mxUoShGYsZq97m5b9291YHGWnaaKjDjkNBLN+H+Bfu8aO
gHIIr/LyUMVjXoDc7WDEFKOB81jammOOsIRlADekaTewN47yzMPWMm49E2KRL+ymPhYcPGlA6QFL
fvswqd7Rh4FUc4Dpz9qmiEIQFnRCl+TNILEAfwSmGFD9I1JSSLmK7Dv5MRjKfwrZTMXRtmCa3wfy
epjonB87xQYzPpQWXa9GdZYFyTFqAOKrZAg5m8TnobGv5FUCJN5ofxTmuI76TOiXkkh02gOC23oi
SDRvqPQJr+6MUP0ZArA1fE++ivPfwXUCcjIS7BRxktaS93xEI6o5HJCpodJG8JBeyYfCGoCgpGas
1rcdQcun21g1ksR78uAL8h+SIaIHtSrGftUvQwIHrOsXJ5dqteF/4PxOr+pyBsphh+j+ey1S/7zz
0YhPFowOkp8Fa+gvpY57r8zSHFViQpBHanxUbFTFDZ4BSPsxlSiLSjfR5QGhhKVcd5qokQBwGqxt
DleyZKJRBsVBklrniSpBWyvdRxWjhh2sDx/RHjHc7YdFKHl8yE+SlVFHScg+BXgpC4sj42cYg2HE
9WlynRZXJJ/JXIQ9iT2B3Pet4XDzkeApryXYjIYg0QBBG2QPqdzviih7YPAvOQ4lv3FldFPxEFuA
jujb89FmurGfp1ynLFl68bo/gcsU1ITkIRcgggb1tb15MoNbavAF5CmKbcucirwMExA958LWP/xR
OWKBDSUZKNsfao6I9wIjO7slxY03472cShL//VsqhoA31sQJ7DB4nj9nIfIDfIu523DO0MLpLYvW
heVFQDQgJ8k+fUL/yV0v1+YEh9epKTrbv5rPkX5kGvGwzHmlWSK5kYmDx5gR5stj5ng8IqubLUt+
X1BUu5bBbq+mOCgQiHzqQuonB7Z4Ff94q/4eLq+CzfhV3lq+6AcW0UclSUdAEV1M8j6SNUpQYTCf
zeN1NvlmQnHuiSOUzQV1RzcrXZtqfK6lxHoKDrIjQotcOP4OJ1HURR9X1/vTtkR5uJ/pIP1NTAet
zLZShK/u0DVjr/R0dRCGgMQZM/VBTB7JSww2ks+zUDBaroLxHS49CNETx1shNOstVx5+UH16Ftcb
wmbEzyLTmma1wAnqsQeBY/Qdccg3UddvVk6IYiiCEnG/mGOTtBZfvF2w6Az4S7926vWyLLfCKO4K
FwRT+lG77jOxLkeXqTlSnUscuITU+wq1/tSrDnaoCAIur9KuXg+jRkw+kmGzlWjo3/nmf9hos46O
zv3nz73wgSwk6/vjZopklfYZCjeK3/B//5HolEQ8UhrFo1a8omJqkSeTySN+zS+68kGey/4CWv3O
urrAYLj1Cs0EQYTEXYvv7cKmYIst5Li74yhWhMctb1HMC97tVAcbdQ4aVNoUWh1KKd+ciU+gS9YB
gjr5oeS+z9hdDAYGnZC0Su3fPFthN+nAfwDM+2FF8+MkKXrvX786okWyU85YFvR9MRKkVWMLxSBM
WdbQtEwYG5qJfQel3Pk6J2bI9tviemIphCMlFHGPdLxedpi7+tUCcPVKgbQ/bVPum97pvj3hpWa6
oEDOdWv9bpfusnT31BWK3LOLBz1VOpwaNkbGPwRDfkLnNING80J4a/gjBPiqhcJfaHcFHjj//bPK
DCYCXOlQ7mAKVuRVb2gUExW34rAjoTtA8A+0EIP4qRXmocbSBW6g2kZYg4whGmD9ev7tuXNnNF8K
04Z5HLBYtpkbKHWkBdyoA3cu4J0a1Ms1aCMlNzE9UNifCVObV3JcyeTnW0GB/AHQ7PlVdXF6Ecj/
f6KbYkTFSpoujNJWasJ+e7CfzwGlswymdVqe+O85OlIutZNIigbYEkQOFHvPR2uJIiHMO18VVoi6
p5gBn5VIHS7uUD3iModXbdeSfiGc9s8M6IlUWlH9czsVRSPFXJjQ+YpXgsMCosTDqx9m7z5QJXYT
mzN7RDCTWVHf2Mja0i9kxUgkqVGJ6RD182I2eUsO5gqO+jHDKAit2UlFcoq5saemQ2TtGimGBkKR
HqSOPzinUUWGOvdY6yy78GVdDk3uuf3SqD/DXs8Jd5TlqylYHgvbGQem6DZ35HN2EQ1ND817gegc
sGEUZ9cWP7cdxR56BvhHbDLfbL11dZhnmjOmxrnQlCitqPWRVafFVkksfcBNrqZ4tVCElZ8qfg/O
fet0hRwX9+kDXsimRIpXpgXcF7s4Z+xZBzlaOHCLANuu9/Tse7cImYLT7EUwaKegtLpRDyP5kdnd
p4wxrdyHB0RCyKKMMnjfL2Wm0XZqnM8IXfBkuDri11nLpuDNAgQMlBlEUBJs6OOb5Cjc+/zdAmGX
OzNShVD2eu0XERvtN9P3yeFNpcRaCzN4MnSaPn64XLotpFp9+0BWcJVnD/vhy6SQlPCTHKUnQ8no
0bbjucydbca+mP3oyt03AqSpjY4uYY0bTf5y+v4KlJdDbUQLYrZ7/tl7UdzUQYTq85izgduC5QDf
AzkaE5nYsaapCuvr6NGP88qI6smhI7SubPohjbjUeMlikvmDq3ATW+HGFRJadbf+9He8UVWKfvxl
CaDa+8RUuLvQBT8ZbvN0MsoQUJ0BAL2fHElmUx27ZyivRZGHBGdS+WNtxJ1sjAxe9jsRzRwi2YW2
+o/QgWMrFeKW6EFnNR+nANCyaIRGeBnFxgD9JjWA1jeoC41OSlkkVNtNK4DHP1WYKtrEAL5jxAlc
51jAe/EF9n1lQGmesc8MhmvXTvIxi8LBaaIuN3mlkXKSIkS8+/h1LLyOOdDXiqtf6hGPAyEBz8Ks
VpDZjRg2EAwFku5u1aqiv2ggxaLCCihgrSvzfPNNv04z2jxO+Jqzd5WYnynvRZyyiMftevkaAAJc
f1leJvsV1vS5uMH7gjnZMBtclzntjZuxd7XID+ZGlyFSF/VENOoAAytCBo2V8rp4bt11W8tO+GIC
gqH72bahIgDETpv0SPZBUv3LvOAa5b4KCLyI5nlPe4EP/nSzAeG+d44j/+tnkSY7K2UySZ9nMbFl
rGs6YnZvgetsyrUyYIoJglalw/ITd3/903NruKSWxoJ4bVByTRiucYwuj4VZyctwUONZKIfLfzJo
5GtfwOteRoCdU2y7qGQ9dasERmXn7f/KYhgF4tcxLU4VURlr2KL8dX5TnwjEBmJ3dGhGGndXxWOX
6hi431IZPsg/FgdjX+rK85n4KfT7FjGH8ukZx5GRC9oQJqGrDCHf133jLaE6QljUsB2sZSy1/LI6
PzaVJHNLGFP8KZ3TWEUgcmSVbudRQSTAM6T4xwGCBR+VgRguu6s1BfdVF8B6P18M51BuuYoWPTvx
tT8y/lzwBlmrwpmrNTAVAJLAfgMsGTDfYCUI0VwkdjqZRMS9Cxgy24JqQkDiiuQYoosAIh1gw28T
WRcVNi7saapGiqCc8Y7Mzpk9F3NNfX1Wst7RQLKmiFdGETyid7iqPu4jzL6DAn1PpEO5dbkhosaP
sWFZv0Svk9Dw1oScAJgRyJQZt/AGjtaEQsCNJnI9aDh5dm9NzEAV9BCMhHBpG2sI8uLGCG3nd15E
Q5mDIetdn4m7u8ATwxpGrmdVYATsOhjWOOL02basZrvgAnrl2RVDM5RKWRaZV+s+TDlcdyd70sFn
NwSTUvjx4XadyjVmHN2oL7ld5YlkBcz5E0IlsitRByVD1GS2hXkt1KhmV0yu62kID989XYbtFQgR
NA5O3baPAancoxOKrcBWCXiE8wKo+gGfV2FpBE6XqYc6OUIQuT3jeXGW8h1Ku5jnWQVCek3/0A84
PgFquglBcoDzFWmIrJx6uC/yEN8orx/htGhF1zI9comE3T1EZcQNM2w5+1WlwSof1z+P/ou0KFp3
PTd8R7vVkV37vRDEoKWEBOs7b3Jf1GdkTNh1LEy8ybw78A9M8yzzbBhtpRDU2qNHxHKMoPKHjKOz
0UuKIaADu4fIGNUWV5jb9Ox6Vhs475PbegzoxaE+D9kGsF/c5IfoXrO8q6o9orsvDiuG0xu3Qxp3
73sQveEjW/SPeAFGThH0ThO/pECkwudlxPznaJjJOhE/Q8MLFglX15tVUdVAgfbjyceJ2RXhyeXQ
7Jqt0NSm6DmFhmE9aVP3GYt3qHamDIdrlBuSSVMpChpV5bI3AkKPIpis790/q7/uLKFr/9E6S7SE
BoPaRtxRYnUGlq1kE2VVpf7ozgQ3j/R1f0m7G42juYh6Nqdd+uypztUZ+Kl6S0W9+F6sPb8ujZNL
IZQUvz9waFn+XaxT2B1ENJWEXBVyr3mCOiti8oy1ncYAe5UDyd5TYJN5WOKL/tcbuGtGnfPMxxg8
aYomSiyKgPHJJyTneaFgJ+5GcG3ZUazqT85tMKzQUKegTHfTgDU0SHGvTSob/yn+URpN7r4giarI
EuOxmD2x2YYT4mlVxwRGJVCpznUSAO4I/lpPoubB3OXJIAzjf04pA3A94dNLznkDVyy5KHlAN29K
990uGoSHugqpEzyCayouAgCwb5C78JoFt4cfcWp9mnDCwv4OxJJeAA5QTFMuLmkmIAM83NWYwL9a
OyhlONohD6pw7b702rutyqRrkmA49vq5TXsjVVELhgNNHsDbu5YGSwKqsH90BcNUkQHtjiXTzUmR
jVmntQp7CTZtrBJrbndwM86spLnAMIJcvwdTRGXvU7hu+tYTqLILcKWEDW9d6iGobl9MS/BOOmuG
0jOGeuAKiSJmjWwthqjmuUPgMVGqcJZ+aB0csRVcCeEbKJddVdfuLzAhoQ4Xl4JAeHPJKV+JloS1
Iwed3cERP9vh5NM8oyOa0+UdZ/XDe2tepCtwThFioswByypVNxzTW8pWjgXjSOXfLV7SaUPLFaFQ
svH9efZIwKUMQnCakJboKX3PAn+i4iMZJpKZkoxw7/WecsqSvmGHwWs0SKzP5+5MSdNGxt0NMqQd
WREKATb6Ey/nex0iSNyn/atifaiv606XvR+4e83nLJNEenkOJA5X+gAb5WLl76UKUm/MekWFr9Qt
NeEbTF7YR8Kj7amRR6vDjxU7+wRSY8UCFC/eB6pLgWTzamLdxxvQ3BLAihCPh7PjPMzEq3elWI6m
nZSEh5mzlXw0CG4/oaBKDbumWOtvFzLrhTlnx3sHoF78/k031twBiLV0ckQyi+U0eBOHXwQt19N5
VmKR8Zz3meZ3l+prgafBly9n8nLTQdDgiedyxRBUA6mXXWu9umAKgBnf6ZHoBi+DdCTx4bmjaiOm
cqmTf1wn1S/NKUjkFRTanXbr7MePKHI+nYKfWFMnjnKC9j6NIZinhzACnor+lUKXOgCo3ELtXURM
ZQ/78SNXXEOnU4CYBxKW/J7NpAwKUACU1WbDV4j59X18noYzWXN85cUlVM5KO09DYf+ycQtKu3Kp
5AYvljeHdo/phjAVdX+OW382SQseOJ4OtZcfGdE+fsWKYO1UjoI0YpQahFoFlF9ObQPJvrwq0CXT
pjrs2oY5GOo497zR94MMLEuP4AxD6Oz3UJeWd0UdyBwbmIXX+WcbKexCv5Nv7ztZoXCr+fturaga
psITqpp60iuxT34va5Dfz4Z+p5Dwj9/yfwRLlPnb/4chgVOKv6BZY+QwBHjF3c6Y87NpnZYtfObW
Tz98RV9k4XgwIxnErMPVPcQvCGI1pqCQQxHSEfH/xReeHEnvX6ZgwmRop3Jb/g1NJbl2lAObraPZ
OQF6fm+NDtZxi+V+Xs+L6sl6HpsOD+/3kTFshhVeTxk87e0c8yJq04qA6gUczemrH+ish1tioaOi
ZT7a0UqkB3nnoRTgvry2cQ0q0omiIXqSezm3ieKpKCXHKRqubYozE0zkTAyhtGQxpvIeXjO4v0bv
u5BfDMAXz4PT7Wuux2Gc1xUi5hp3HDUxtcT/+oAB3FpBXoy4NXtBFrTNFgaHEMkJYM7AQoNx9TjV
NNWJamSx1aJ8Alajl+lXKQBdWlkHxo+/zbkdjaIkEuqqfTg4uXG8dunLpsVVRU5ebNn8eJUjoSLk
gIFcU/j6+cVh0yU+l/P4yYZ41+y2ZRknRH5PSijUAC86A8VE0Uim1exg1fF7iPm+WGvPcip90/Wk
17lvVBVt81BGpFLKsLp8WpbMt1cAsjZD8fa+iMQC0d/nsDwRwS2aEbdOSckMaJEHw+lX0hcxd/jq
bDcNPhZq8FUz9wc+vboJt7EvizpZLM4694EDGYxw8mkrZw8xTRxIA8LZeJ9+hgKghAanXh51Q3PY
8QYYOrjCRyFQj5ksFHa8AoeHvsbUJcu2fji1pl+36PS8AE6ctUS+it26ruF8b8tHDCW9YhI19gPi
jz9979eEyXb7DbH3kKBs6wQM5YDpiJkXPFa74DwXeKTzK5k7C2out2WWcFDgyj0zLKu10xdqG1GG
yfLvYJWDsgsyyNhSARnF/QtyD+XDL11DbPCDzsGDbA8vrfD6WRl59QY0AUbZPsn1nB639Dd+NQrv
IqFDSYrK3wFw/2lOUAGqgnK4t3CKhnXk/x20AxRS2Voo4QlTYwUzsuOdUlH/7IoAMOybgXaApMMb
3y4AA/yVVCccxd4/VGIQ48hW6v3lC1XLqPDjmzILlF7eFazeeoLthGGEl2DoxHigfVhVgzvh81r5
/dwISxgCQkWrq3UWaJXIaCz+5M5VNo20OJ7dlBNYhwEumxx5rGW83hIrbwUVxNmfhSzqpB7JLnL/
+Q1cWhE8cgXCtu5jOp96hDunRzVCvmGCUxWTQpXbfmUbz30aRoIQ+8Bz0NUZxaRKYY1oao8GAVAi
DxP7ozg+iXqqJFnJdXhHamIjG7mpaqpVnw4i202XE9HVq/CB+YuEx0+AHFc1ev+tJpWX79dT6kXO
KCTT2JvuWtQcNAy+tcgFMMJjltO/Et03ZTc4Hjz2lX+Ryk1RILbJa2KRR3bKggoBGiLCBmAesDoX
+W5s7AFX93WdVHONACM5EhV76QD+BUJS4BKcsa+3S9A8nHlAKqPVZC0uDFmEMItoJmBEFvPTVIwj
Waq5V0VlCxD2Jbn7syVhE1Og/Iz8u85LN2OIHOZoZ4u8BFN94RimGse6xiAJY4zrGjgJjUFZhcAX
ThlXt6FnCTlYNs6NVjFTQvZbamt92/xYe/vMP88z1RdAo7ZuYhLJnbXY4lG/fxLsYdZnvbmFvT7L
k34ZPHmf2NDtKgLheoS2F9zkBWPO6d3sOzb75dD2cgDoMPwG+IaKKnPcKmpybzsK9ui2weUsR6g1
bsvnQJwIfjpPVAi0/38YL/nR9hP4Hz+nHfIjvfdSkH007QboKM1gCcLKiIQvZNTxkWXp1sFp4oHB
kIylYKCeADVcAG+97ZJ5T9iwmU1q9HINa24G0yKW/WzCH7f+wpKJL5O9dkXt9p8P9Gtbiyx2sG00
KoowFMyylyqaL0DFAr33vn90KsXlSYgoWeJGDICZqVsQpQ9FFlW8kJGIcdOHR5Z3RBAzwuFxzbse
DNvEiOU8XI+9joYByCQfLGXPbE9RZPIAyE1mDnCDb7+SZ5rtsN8kmGZYON5ZyJKBqql831icYEZH
uTItxzCu1cpcGVKpdUaqAF/hRtfI8PdL6DpslTc3QGk8Bv8a2gU6HBrqqrdMpspGHbfSBxp9uvR4
Yt/X47E3PISDThD4biFum3pnyqnVtOH43kB0QoBPkKbQkM28PS3RnMnGgimKLvmF6aTO8Ph0cRIj
4ibYIyO1mmnWYV8fXEjTubAwBYL0LgqB44Dwnxp0MgMqB7Sy1hOHKC0mM8BfgxvS3BKY13LqucWR
5aB4KEIJupGDgKKUt8woEHQKXMicpli5MBGAp8QMF3nAMLHwRmdzaBTCJu2iG98XLHcWGjlPlbj8
fbMeL0hwbt3QXzoyFrpIslkA4V0tKLPSZvIuE2Tj0q2NXd0waZT2yebhpuDXQSdbdKrWc8ecG9Tm
epLcVRjNCtRD5wO4B0SxfArYQL1oNjqgQjXsk99zj6yWSHW20qGQYu08aTmVyNeWrEbGOZqZzYIB
pp6F7E3GTPBv2JzqRmZM+Me+/2+5hMILIU+IPeC11sLQPUsR4rUdwP4upvAZuFAgkKZz5Czi+9yM
m0vegxgQF77+4YeY+ElDqzcSJLGEjsILAV1bD8i8EKX93IMXtqjj7tf2uI/fabt+uIhSc0md6zKg
DwOcws9hOLcqL4zyEokYDDVuAYuqPiepPeXAeXvFVvJeenkz43RmKZClxEKUZZdJT/R+FkqgVVsD
2zSayH4+mF4S37X180FW68KBu/7hMg3U82nP+FPBDOUktN3cwFu98dAGCZebVYfdGkMXTFgV5co1
tqLYK+G+dfzFSFMlCm5Ofd7ODub6YpaiPFvmRG0zY8A6hIOM0fPkkVAet2YA2Mb5ZCUDXMZLUQJ8
fWa1I+xJMkeD8HP9GFk8kbpw8hyPXlC5WXlmPQbBVkCWaCXxvXPJOTtYs6BZVQwSsHcuAp+HJNZ5
FfByvpOELMW4BlWwMy4ypZaN6+LtyjeTGRibgbYMRiKNFGV1SXqwpmgSlF2Ar/3dd5dhIro+7QrC
SQXPUvRU9y3KVzsaX5uLzxvpkKlU3lpxJ+vaSATkzYUn4ThUEl/8OxQOFP4Q846nDzqxMpXGpnVs
yCGRdSIkcqE3KQD++LYN+MrRfDURVX44w9lhjbbgsumDe/ArzpCv6AjpW8VLOyDRXCfccbrD2Wae
6GsNcCdkL4llcs2wELeOnqOK2K3Pu+zjjc66FvYRMSp9FKqJ2bZoJ5p99+JG7mFOvbNk+14HHt2D
ra6Tiq1k4sOG8uJVvd4ZCAnVin8RAihIFr+VcI9nlz0Itz+zt4lzRmHRACqeCV+KBzqnPvXVlTGS
L5VWAXzUCnmv9oqAVJaWmV1JRwbBNH8CfG+qtGch2YVp0rlDDRk0ToAosJWpzbnNnsllKJk23vv3
lwb304hhl66hAbFVTijCgC2vIEjW/J/nYoogdWghCC5791iF3gQgF3O+pTd2mCmA+vMH79kazdMv
jJ3xL6LFboOx7H9hQObnmBIhgphyD3lzmCxH9rgGX91IarFLN962HfDs7WpG0zsN6sQwCvF7B85+
VUOP57FhusOekydCCc1JlqiIMvlsxzN79ksio/cakWYQF85BTGPy282qR1eXU7NsXlD02ao+lynA
5dRbT2TDtso2vLqwfbt+GMBJ5ASlFPT8uZxY8fdAs/hH96Bi4PRyYv3Q9JTLKGLrxHCHZtjz7lVu
VO04+5qOXoNMiWExCbQSqYLxWVk33tGziaQsgKv8SU5Hu8IynZYaB0RFgFs6OjY9I41C3OKPX8FU
Md/zEQXTaM629TnM6lDSgA4AtQzRljJmv5mwFu9jxLN4N/yWf+E5co/jDcBaRPz/Kfq0Szt45uZ8
BajtUVRVvjAw3XFh9ZykcDEDPSzJvVqFokK1ol39TN3FTr1bRtWdv62iSo9T75ZbkY1IUp4DVb2n
x8eUADJNfCJ70aZtk49EOAPofiR4rfV6qliwHFUHpP1sS/o5KAtBKD9QyzsntXzkKlCI5FMz2s9m
SjGkpuJ4cy/7WQ5rECGNYBQq31P1SzLhj/tU6YkL6YDHoweb74e3qgPRWU60Jlv7uX1Tbzzfsv3L
Hilbq9OwNcWJ01M69dZvixO6U+YDoQ10nizQ7kxJXj8vLbl5nCOK+pruJ5i2F3uf+QSq2+46R2XZ
rXSBQ/Ti3o9chTFbYNIcrjpfC1vdb9zCG0LsG0jxk4qPT/glYCeIZ4htD8CI3ba6wtQH9eQKB82K
fftNSKxDcR/aFl95CgBrncGCappsF1G8tjz28s0xtCVDBSNpoIm1mpMAMu5mzJi6u/6S/AcsHMc3
DZ3v289PDTXtq8NsUSpvLQKZgNtc5S1+QibawMKQpk34PmpPYXlLMmvJqFWTbo+L9n+m3+cGudvh
iVr6GXnEDOOnOu5Y9quMU9c5SGJVMmi4BVFoB/TLYP4aZ+AAWSjS1+BUHKCg+e3cEV6qcBeq04zM
fc+KGK5LaEx3wCioyN0nT81PaRPpcTQGYhvXxMV0cUu71OqkcnRZ2M/UodvEqVjCNh148kySL3Jo
BS08VdqEg9sNWh4llynKf7MkgHYB3FOWfnDI90cy7kLMGe5ICk3RU8Cbszu67dGLS92JNHr8KrnU
45e7litVHnCH70oMgY6M/Ho3CVJifWLAUJcJXzzdSl2g69R9i0/UEUMLm3Rn4fXzwwqteq4yZLl4
9ayg52MquQH5h1TdLubiNOQlhKgw+EQo7S/EjJ/VwFBfpuCJOezna1Y3ZpG/vXOQnqyiRAG1EQDE
3odDMNHWW1WhyuXzdBLJr5nXaa+4QmN1zm/3/34iJykmXu2WZj9eDImHMAIhLOIloyEU5w2F6Hg0
vmJWiiCKaV0WphJjnti7yF0vOQxPXDmiVVbbuEnTvKyWooFisIoYC/bBhjXWak3OBXtze96Z1jKq
ABUWlO+3abWqcauMBKaABQufqNLUHfFlrOaMVdoosCRO7LH0Niuk+hfx5Y6bmyD2rQdSOwb/et7Q
HGlcgEXlirGWbr88odWiT4mglnhp86GOtae/b7aGQdc1fOrzLGcc4QP5KpowZaoum9w5jmON8VRD
F71+w8CyYmToifXgMoE/yrYq7SwutsqZwJ38ihAQsIOV5xi/fdVMHS7RuU0aoYStbtnF6HNyVYRw
Q+ttNN9kFkf+9BRaaNG0CWTKM6oK5CL8Zpq1HNLexvILB6CDZXvr3TBz2V8+hhE1MY6sF3ZtzDaT
OKhEvnOUIDPfjxJ1+TICYwy2HM2QoGiBWYC6teWoosIELenjgZkoq0GB44SsukYkarlRZNwVtkYb
p/tyu1gwaEOPwtKdaydF8eCdkYd/UgQz3oshfbwz6v/gJlvB1oDSILziJFaJ0AiSQxGntr0FrVDA
drfZ/B+pxooGB2nx8TJXqeaRlf0igjpGUREwbhGcITRGm/yiieg6heucBj5Qh8oqZWBME3JeYEhl
Qmg/5D3g+kAbTrjyE3dekdAt8TcWe8boLBdKIX+cNbKpeUDtKINDLp9WNRYYZFsteCpzKLBU0zXV
pbE1T7iRj7KixoDj7u97xZR9QWqhGrpTjtCD3a86RFyw5oPpW65iYnMNpCs5P9JbESDYpjVGUKEz
1AIfKS+Gvj21zVxxHRAtMebxso9PfJSRXC26Tqxwy6y8WLPS/POehGLTxfX726f67JmVaBnOriKQ
cZTr55cnBhChJUDdafdRKYfyjl0iZ0plcvOe1fsAKFq1XSErD/d/C3erMP/OrDVwwV9WOtNJzquP
v+9JNOTr3Ab+WrsJuDmAQuPlqHS3Pha2YW9r8eJLl9h8Eq/9Hl70sX8nsJFtZpCE220SzeNCEjX3
UcB7/dPGafH1YyPIGutY9lhAIcMrAIHHXSHk5IsSh/QhqzB86/mRRPhHqp4e7bikwU0FwC/YrCMz
jOSDbROqPhzcmVd0/n5BykKjGlHUCr29xfIc0WxPRHr1VOk6aeLAWHA5zwkgeOE+SKoF9XLj7H/g
cYMH7R6ZKmXGZGTg2dL8pSgRMdAFlD+A0F38TCT+2c4IAUZ1EpxyA9PFe0LyGhpFvW8kpJex6q5d
5h3DBWYZXQKGjG3SVnnRVMDJg+cP7AcMCLoIHMPh/ikk9p2dVA8zExfu9QwvCT5rTDUtHYeZhWlj
6FryUOU/Pgz+NopQO9kkXNXkv5rDiWsHlS0ka96JyvKehYC0Jjf9T6IMJPjT0kouzim3cyomAjns
C3lIar5z+wt00AQfzw6Ox8y7Tvj3Kxpk5xay/uRLjLOxmrE97fFFuNOSLcFDPtiLbxhZCO/hj/xe
MXZOdrcAuXjpfOT9Xr8kRoBeAz4maSw0xAJodQwht9wOh4douHts1B0y4aqkvWmYy4mTyBkRrchF
LSp5CA2pvKlUSoPWAktx66TORJbJI8OEgCyoP1r7s9iWvCFhLZhkxTipW3yavoVHKRpJKnE5v/JA
lyE6LjuDxuFilJPPikOvN+rcRFJQGeRfE9s9cKhAcFQWTzohTdZ1CCQGkF8Er+jiXJIwF+Zy1LR/
cAXmYlJEc+MDLVVMt1qwQEjxINag0ZTjrJtKlp5VspRa/SQtLQK8bH5fbk8R8oLnvmIuQKF8WggR
F9ddYj4X2kf685zj33gP6Q5PYGL4jABC87XdFIT28XZfVr/81/dvH+ShKy7Dwo/qntx2g+xvTtZp
B1snYZFQV66r2M7O4d7KyolpKWEld2KKiKEg1VQCsHCTtR+rTTmfD8A9knBLGfaTFuFVg+TOpkWg
sLUTvjH3c1SzI/yLLS+gCc9M+4h++2V/P9CGkWM/pC4RxahuidAIzVrHD7iVxMfSwuC5oCrMUFLl
gGwMbFUbjUb/DNTqS/DJcggVgYSInwsMyB2DTwWJuNin7jBVFBf1vMv9K2FGBiLl1Gnf4uogA8xI
56viVTfsMC5Fum5Fr/7A1Nzwsu/qlWuQGUXtEDE+e8wlWPqvPy6xgzmT238D0Z8gDOlMCr/YKmjv
sJ5T09wON0m60iBj8GbZRQ2q0ekpqFpL5IxqUIiXsAqxWL6COV1kpA4IuyMy0nNB6P74Bse1ZnNj
F4ylHxrOfAdCZ639G9d7W2fR6iVCP/c4UB663tuSd2YTqwXnOTKKEQt3KmqM93cXmlNNJbm1CLkX
eeC5TGUGOKu3mBDBTqp6PLe36oODu6LBnc8EPuGpOr8n4aUy8S357AbGm0hyTuOBJFCx+6GK3j7Z
6LX3rp6VO+eJiD6ULzO+zjL25fp6vW6KvnNuMn0wYilz02hzqbRFH49f7VT3wt+W5nHvbdLf5H7u
/nC2g6fPkGMWbv9CkAD3/U+XkIZksuXYuvfeW9c9IfqKq16dtfYkK6r64SV9RYXuKl2VawrwTj5V
ANgReeVRGMrK/6RPICfjPFbqoPjgEY4t4HNDFN1D2iryClUWSswi3MENz8vo8lt+kIaHyfewteVz
xtW/wBSkJ7Bv2XsNp+T9u3SWjPm8+BF/XV34Fg4ertcWKzLBE8U1435Vj+l/ct2MikGGqKZ5OXLJ
TlcPzQrqK+fOpoplHYzdPQ4sBzAIOY77AepmHc04auAABeBohZimSdgA2MwOrIa52qRe+xunBdWB
Mbbo8TXNriwaGf1olRyGQYVWZEe6g66Hor0huSPVZqgB1/2YR1RvETcEV+Xk/ZC9LSGfsJxSmztQ
9IIadgApNgEOV2JVV0+SriRk0VwvryUcVtZk/WQBPWLP5Ykwod2K5kopkWVeIYYs2CCheim6ZCdm
TcGsuP9VzJlSJ2v5jvhMvxT8qHQdnYYtC/1Zsc70yOOZJkA1fRn1MNhn83wtOOUdvv0CWBwRsJuT
rNS1fxWmrVvrN/MYubySviWM+HlZOHu9+OONL/KCTQnbRBZ8I+n57tebsKEXmi0ZGuJf/MRN4v14
wMOJUNpZcGouzzlJhNrhpGjrOVejWGQWe+XV6SEdcODwdy2je0sDtUHlE+kYjRPEoiLST+8dvfsr
tVyueHpKCfU18SSWpzz7nbSOyz8ggvBHnwaIYwK0rRPEbtnB1GRcMWL7vVYwSr5mrIqTN5BvFfjk
M/ggHa4CeQ/2T3/LVoS4SbD4N73Ihg2yCKl7XS5eoRZcNXyTgyA6bGC8yicjpf8NobOTBkAe+PDZ
SYEqvMFACMtSuhMi4WxQuQIYqXCwlRDexVXiO9thrwueBTRcebWLa2nYEKq/JQPs53vKB/QeJcaf
IxENOThe/nwDyovUtgD7opiHKC/2hAZAUUrquK1CC+dD907iHgZXkQh3AfUiAGW2JbV52A6Yo1CS
NmrZOfQ6Kf0znqrpMPFGJKfPW7QVHF51ZCjTVk+GdYh03ZmEL0KchI8cyFdRl9ra/esYrB7FWvsx
3wsoDn3CrW8Go2OMdAfO1aaFBKEhNOObl4vfVC7NkLOzjb9QCAMC6bW+Y4NcvwxIm3Ni9Lz9Aq+Z
+DKe01ut7doD2kSBwNGxQJbsIFOiqSGNIU1YGK3gAr//IOO2HpEWKEKVZx3z0PwGiaDSLMit7tpP
KFHC48/oPF7ZHoWoesYfAJ7gjp1e8sBqZGYKemrn8ZJcP0o+6P+AUC+S3cz1ynFk61DI2kGNOAAV
ik2oKNo1qnEKCQUBmvGMTKpyTDsEOH5m2qip9fUThQumYzZeqSulwWxxr60WKBMNkIh4HrYixOjc
AReXDCQKMdiQNlvtxXzj6/vhpHvJeHbeewGy/rwzSNBwPxlC5XxJPEKPSZ9YA/J4H9rE5iDE0dOd
lKhcHPqVUEwKAix05lokd9IHbPHzxJ/ap+9suTG4o3KO4o+RHiVmcXUBPRAf2+NfwYhdA72Bc2ch
6a4sO9w8cv49/JavYX7Q/wCj3FuXIWSk64Hn3g+qffWexPX25zQSpRH9rc52vy3pLZtpLhX5uZJ2
EjATE7MnC5vVomw3O7IfvcBnfUEUdL+XgBqq2hFnNzmxsE0XFTiJ6kRpOTx3Dn/MY4Xpq/hf3m5w
3c0U/2NNPAJzksNOqPooYLnU7Rh8QZQG1pANdEalWA69v/uq0DSWAl7bFF8pLUuSnCdN7ayJlOZW
I9ggX8/CENek/4hFWK71dMMTRArsKsPSwqlHphz+bwiIu1UsQbzUz5ffZsDyLROtf2N0r4s6qCTN
aLIALtEDipqWKYcnL7vsWvw7nk55h0PdN9L1kibjRJLxvak4Oj2LkbniYIYdpaYk2af1H435eucO
yUhPf6ebrs9ZFBFu8pjKGMcknGbloWq47NmBrXNRG5HLAUT3g8/Jz63PCZZF4DmFbr4GFB+600oO
HTZXWpm7iFXd4lysoa/Bz7eogmeWtYCKgiWAOfHdUqDqHeptMWJ/H/Y3d2OyaSozx7ECYEx+QJQj
tvyFcd1ey8/hI1B5A8yXwjc1U29D5iD8edS9fgwGE5n3TtL/x96yYnwRhFR+k1Gyjit7I/ygaj/R
Ud9dbduZ00NXJ0nfNiiedhuaZ6nCEQzXBznW28geBUJfLQCLDZt96TdlaA4OCsX0G76lVREuOql7
xW9KQ/wezZK5mT8FcRfPwlng0zQmlxveycSxajmf2b7mAunWDBZX+ESv0KXqE8BhVsw5Ahe33d2N
DyTklimLZ43KfVMKEIBz2COv5T4poGLGIIL0QzMV0ItKP0qYzMK/of+/VDRmvqEIXrjpvphY1aG9
K93A6QzkTM3WUIZ5vxDT/R5ub1c7gaqxFODhjeLO6em5W0ScYzdVWapQ31Gspf/9XEdEoIHb8A1C
aW3LNCpXzWl0jSsa4EdWNhKKlZitz/LzDMpJcaBaObCmT9EZ0+7nWSkFVJhV9juBfZepQsm+tcvn
fVW7WCX76vykB3uMCaK1cRjRGaWwzc+CAJ0aIWHVK+wdEyT8SyaRqzp2zf+dZSqbwf4hKH2ERiJ6
2Goe0dCFgmhOJyJnhI2Debnlfu6DfodjeOGsZzG94moknIWg2aJwaqjhWzFpfoybbUA+lLtPQNAs
sjtSHArL2yf8y5Ec3agQPGYtQ946Pm+4/dVYIbra2KLIJ5LIcLH062fMYU5Tzo+Ygoe0HnIipMg5
0tvgMu6EBRQ23Q3JPy7W6HFPHSUahxZagoSAKUbVguXXX3J/1PVBy1ltPcBc1fneimG+iWBCqsc2
9DW0z6xdmM7CfUYLb/iCSRCPAjybb4GyiPeiYVVwbbgV2zqyiWgBpx2dBlww35u7EF4g8PHZFaO3
LVUkACbeqUS0qEHEHsREefVSMsRRgBF37xNKNM5sBulLwm6GSkX0AN2zy9ZmvQZaiIjsnWBkzGLi
sJ5ZXduWYLMQaKkJsv7QyNGbrrt5aKl4HHeofIz/WE1FMl/WIcnfyNejlDH5lukc1a4mkKGVDVYL
Ew7Jge+rKJ2eZPDuzAvhJ4RwwW74vwJFRqAjmxpHCWV+/zmdM6f/JgIQH8Un312ybFfj1VOkZZs9
Bb9Au8QWmgvzNxx3QfrQcoj37iN92w7yYN2t6hZdczhNq5Svjm8gUfiXsLX7gdF0Ve8sIvzLyb0s
w0VYdTN3rMRaqxYezW+EW78j+PEqQbNsnckBw8aXlK0uZ3O0E40yl4pVD7NAkYBZ/xpFp+roNFoS
9RuWMtxcYMuoIfE/59z9691w16cPnVtokJNc/AJ/ka8wRmXWynTli4UztS0WROG3NIXO+5z3Z2xB
0s9lqiHuWH6iUifddGXryTqQpTWg1tNL0sYi/FSPrqlEm23jM7vS2riE26lBuXme+yyyimifPZw9
w/3l/p/yAd3bNAzOrFLBlmnBQB76uKiEovXsd/U35FA18u9fYCONasnRYRrUhEpAt985xCX84LpX
3wWSDPmt2qdE6InJIYo68qJT9NUwI4iDHaRoxKRr/mcXuv+vjT8sLKe+Qp/z5Ba0ZSXDK7I/OzrH
OzxG/a8ubFmIbAlUdzjw+WtEPevYEaHfjNce9KvMUn9FfHGyGAD3E9tY7Xn2DxLyfNlOuuaGfhpV
v5Z4k+zOsxoOxhkj7SaQrYgaB8m/+DV23LpzR1Ec0zDiFfdxqsLwfIK3ZLEc1RH4oM2xoYhZ6tES
o28ZdfYwgaPXWjfw3/DdsmXD9DhUvGXurQ1Z7Wusff9FN93gqrTvbZyEkDcwAHN/vQ/3IePJ4Fys
8LHaeoVKAFYFg0O1fXt0yFozVld0ucQNoxtzblW0NMTx4TsnCpPbAx0aLn/ojqLLxWeCjmjwAxGX
9JZb6UoXJEjMoza6YSUCqAqUTMx7NneKqZC+JFehCkNUaGjEEn2Adj+m46tkUoVZ2RuU2WPyPDKn
oihHgwFCXfBTD6qGWJNo+klXKzY26Q8Pd03JrGPWVcysruZUn3k2QRen1277VTmeFMO6xAnRu/LT
W6snoLi93BEy4CFbhwRypJvgXF0KSRvyarLV3vfRTETEq/cpCy252zdZ+hoMQXvsjMWjyV87E6+O
f5tjpizTdMhl1plt7+ZOc+Q92XGXLJmoN+M1UYf3b+wdPF+7bXjZdIS05H92ikfGNz3Cu87UqF4o
CTiRNegCdKWSbkMIoe8ayTR+TLfyLCXCAU5mTMBr+CbRzROHTOxpXkqOVwJXKpRdjeUYjEEwBrtv
So3ZcPzD2p/ep8k1TynA4DVyOedseSK2gwZDRnFI7jm3JpBENI00oj2d8ApkvBk+gbYm0jH6KWcb
sF7W8WJw+5jAqMmvJLbxYdWlv5Rlh9K+76MehtZTQJbC/rdwp6vKhdFTcwPO3Xlxa/7IBmVH5V6c
vDCtq+whlRFu/H4DzbFgKRJr9F9yJPDvy0kB+sMDlsxSltVuTzkxKzzAZ37NlZT+rKOxz14Y0QWU
ZpNdQFeX1GfEBlVsh7vr9IrkvV0hLg9VyioE6oOTWXycHBU6WzIirBq1ZvCwG01VEuUES/z+56n4
jHI4yoPOqIEhRLO9DAxmmnrOgA4Xoo264ZAc0YykPLl4ARDDU9DgULJ1IdoqmiLzo6B/YFwDOWtO
Dj3mwqkA8YtWruSJN6vpMxzmtIbP/mS8DU8v75sgwiSJLDmGhxl7WsYJuGbI4zJQO8rYzs8UXNc5
4Lue0J0WeoyZqPUm2RQw7TPoRCQ4xPDEbWA9jKfE88ATquZh/Nl2jEM5REjLM/Rr3DSD1cTe8SMP
meXUBJwF+AUZki23Q5umG2JKRd/Vioad2UaCaeCl8UKaVv/sX4ZEka/eHfmYhpmtDCS2bSLFS02c
xmWlyq48eOh5ryIpyd4PLaJ1MLSjjRUmH7IsU2IJvZx1k9c0oPiNgAafGbkWRZ7vgohgalScqzL/
hipqe7WksZ/yuasL2Gg2iJuZ9Hg/Qd1U7tFU50BhfTaKm8EZoLmF5NrQkL6ns29+BYxgPog58rze
pRUxgmhOlLZ37AlKNO8GbrAXYdGGAXC6mghqi6teBAFNJZVmkY8bqr6IQyekGMJhYuN7vXFu0UI+
fiJoJu39EFEeaule4CMTlZqvaC5m3+G8LT4tUmPugD1dzbMB0mLQ12RMOrp5b1Fgn0PXjPTm3Bpi
x31K/kxAUWBALu2Xuq93p8G1vbFupb/9YDFMmxks8Au3HUN1CSItrakbi2xh0W40rhyH7wqeboPi
7D7AfpOUcAqfou8n9b20IWxZwH9LxDUANWhPRGS+GdMyXzujo2XFS15h6iUcmMJKmsfODnU5dfql
UeYPVwzKumvLR37Fpu51FJHzDRnasPPURsRdm9a26DPujqxBOK/NspumKwhJ2TYF/7fmyVqi7AKN
dbKuGoTgiVzE0GfRYfDVqYUjOPbzdP1/60BLC08n0wtFiweBzCuFIviSqFZfrpSK0LX89nqATuN7
7YfhS8HQnpiMKIYmJjrvBbOW9MscItrpIV/CrmvtR8ueLt1/rbAIxvunID/Vm+xumZ+zkuLzrcg5
EkqZ78EtY9IH5b21SDexQ/pC0MZlvvUYg2MZkCgk3naXCpNjET5Fm4b20sBJc/O9OhII/LbzPsoJ
4TkcslJTGt4eISxLkqnHfmNZkIf2IUXK5fhFTaRR4VXJvBckjY9knMT8dC8jPsmeireAjTgwG3P1
/YuPJDsHgSb8yXNyjtYrWZLEF7gamBSFxzrVfKkfrQZhACKYIWY8BiTOycEPK9/kB9weasPuHRir
pFD8IcKbMwGiflf/R9K12jPRMYoyoygIEhFgznt3i4d9dMxvgyKEnMmsuEDl3iliSYfWvBwVn1sG
BFCnOHKMe1eiOoX0O43MqGBy8/cFnfswP3dgLvDWkMDkEGNUKNtPK7lHEKOaCQ6F4ehvB1P73ED3
CWkwMZ5Fn/DMLP5xA0hn/7ioL0SYmVarj9722KXMtTn1PhOjBzu67TiLC96i3tn5bFjx3bamrNsI
rfmccMW5CGbIZWvyMyCITkkSGw4PFYxZP7tz5w/yBEjWPGtxA65itLOpnZDx3eUwoJ/cNJl7l6ur
U5a7i/fNutpkLJpyy307b9ux8g79zPpuzmUtJ3ngTN4zfh4woKzkSmKmBoh2+D22pmNLtyozExbf
EEvhYQE3agdQWbmN3SyRlTeTd+OSgqUu1kKxY5cupYAububIn3p5+Ov4l1oPbAauouqh0prKPxbj
4pv9I9zn+Teu9QGV85zaxbjE5G+2X68VC/2fsrMZpuljVQln9+PpVD7+AqzU549R+RmgdYtHV3SJ
y4JcbJTeuDC46lAx+6XnLa/YPnVLB6F9SP7OAI3kgAWBcQ7jVqEqUD450m+vx6+CboWcPFISwmvG
lN5hjgsQw9Em+9r1zYjZOJBy7MONz4K5Bb/J1C0xHopTJvTl/ARHDdLRp5oOBTe+ohVMFtkEDNa8
Sz7VABS7UFClCAU4m9N/AXqPoV/5q31Pe4CkzrpMzBgeuynJn3eIPRMmpy821iW+4GMdP/MjONpz
Xcv6uW5leqhp88Enim/cfm9cS604Ue/elyfpiQRrptAUA17tukGs3QupVw0jn0XdpoaVEam87LX6
Pmyfi2iffXxzZiOFowM1T/Y6zNWZ/k2zXb7La8whWT7a65lgXs+50Av3mdKxNeMjpHqKC8myOj0M
Xf1Hh/cgfErT1tBthj8EB+szccmhIY+XBhUywUim5gFIwJicivr0sOkptbYTP1fSlHw2H2xK17RI
6/QHXIJiDkLkdS0OgXPkG2L1tVvxAqTpapkqDrv06nNq3BwU2LPxxqEp1iDLkHQnB9JRIKqyiOVy
jWC5BPad+Cwv50oL0BmFUsYgvsU0RyhZGOUwnF1abVIYxu16GVet0dULz8vLEFuEfd2OKw9kfBqn
4lh8lXOc3DEoLQGvHVb+5fcFYAvHXfithunibsjcnNYayig+kQzkTgTJcXWGoNoDI5E+JAqarRn/
AeCOg/ZHXjsF/DuD9Y/XZhSMI/C/nEdPab51NAlTjAYiBfVzAMPDBk0NbHhbzvYCXjjgZSUMUH7l
uLP+7ZqHIamhVgyH6BOL25+2pLZ8orcWUD4/Dcwram//EoOFLd3RE9vVEMvRO7Xh8WwuDNLpv1lB
FYnnliLqaXsTYSktZwdeisOvoli6q7tNjZV9x6VyA6e2GpGRWPrtWd4OvoBPqjJnQEUcxY6m4wDq
ck8TZFOL9potMTVTUkjU3ABHS9WkBTT0Ssr7PeMBZhLAM5XBO8cYLa+F/hLRVjuGkW1SlqhgezRs
sdpATR26o+MSR+1OQUyy8Kj0zEjbYkB/yaMathYXOQVyjYNXzgv9p68UmKAjAvjN+jtmuD1uRfuQ
0XGF8IX1z/OqnaEZDpqOGU0go4N04e/oVDkQT7iMVvyzricLxRRUa5axgny4dMi8mgujBzWieTqX
XhpoiN1/jQwInt3+6HQy2U7gYMFitcn6m4IddXHEPf0jfSzovdaI3uhEeotQhqQWnpc0HANQA1eB
j62ia46bR6qTLtk43lDz1JyYeTPMpwbZ2jEGEoj+s43XWUzmtSw/ZwpHT8wX9lHvxu+Szajd6FrL
f3TIs6vdKSaNwsvkTToPmv0JS2fcksUnxji7r1uv2EU7EpuPozWq52RuGLsHwPwclS1VpqX5oqLR
nRWDI+lg7q4tim2v86XykiPZVNtTwy0F7pGBpGxmotEMCO4XCvEVLaJ8VIInKoeROtUKYkUhhVUe
5qMsnfpzk7L7eFLIWzrDv9BzTboIdcq6Y8DzWVhVRtzJUtzexA3L8riODMfRzKAFeTEsSoZyZlap
fnwTbhXvYQF5i1MRVuZxdRv1Oby8iNDbgKEB40xQxPFH2uGNtuoa5TUXeuMgZlIXoL/wwfgP8lDv
MLffOB/0WdiyM17AsOc165Vpfk65hBatLc0Ro9rD1xwOjO8RR/Pcll8R3YFWmc9yeJG92eDMyeM6
7oqTeIvInzPH8QAotusnr3conqMR8Smumj/GJ0dBwyJiwvVYffTTgmiQCVVQAT8BqwWxApaw+yf8
wwVNKQyBnvEvhTQnFHM3uJ7XdC2FeMuW9oq/1OR+qkdeRd8I8rAuUAclR1/6B9VDu2G/ZoTmLLGH
adEh0UgDRtBQbtFc58Laah/6of1fECM+8Bia4J3sYlNC+xNm7Y70u1htrGFRD7krV1bLXsfaTsWR
Iljr9uhWPec8kX1XsJ8bv4wWl0gIpzb5edv2sLcWHD31pg5K4g6/4y8TLhxFEkGVUPKp2w7a0j56
waU+Y2aT1hkb4L8FM6w/DVM0HB6N3/TCSocBShUCeDba7PuOX443AeUiSc1dgXvuo5atzsamz76o
g72Yqs+ljHHqbiFfvBL++n0ApwqG1EBzyVyPFfRWrFFc/DjZfWfvZDAmvzDQ2Cj6IqWRmydjyxUy
3u1XDnV06MuzHJwRqZBP+PXxW+LU1z3ps1zAcInD6UtPhwm9IV+fC3KO7YlpsoTVPNnQ4wtgVRww
BRTdOU60eVZqukDy9KQCgsqCxptfhNrxOcpAmKsYIOGt5FztKNe9+yrp3AmQsUpSgXn36BVjHoo9
Pit4eYcuu3+JU6JI5e4luEz81/FDZK5/ynMvYrOBdXIP5W4DPA/LwvDJYdT75Pe3iiPxzktD6++f
7xydnsDXBlaj9wkQp0jDAMc4OMpV7IYKjmu/9BI0C8mE13mfC5MMl34bNlZT9We+cEF4XkWJr8Q0
XCu709WJ41Zmbo9Du4W4oQ5cyhS88VSoexF1EV0JGUeEBvG2WbECapTF5SHxRK4LrlS6nAaeUWQ6
rpW4FdKJiH+NwuP+LCAppbicrK4SK1/L/2jTaFveasGSoN7ZxEzgHYXDl2Wm5lGEBHrx8ra3fJqt
DSb57e+6vegWg+3igwqSMiShkhEMGIfz2c1R/QFIupQI8Xmw0tg6gR4N+POT48WUFS8LaJajM/ue
TvQY/6rA/3pVnn6NA+GC1UKimJjMhb66ld91qabLTS4yJSKHdYBDK1r/Q7EUMOUIMwToGkF+Qjfj
LbqKVqjxON/UtCzFCnLUG5XYzKRqo6ONPHMrgrOtIHkuf93EwTMYq8nHhvSoWUt//AHvrKcQU1xT
lFUOf35VjfRd9HM6sdoMQ3dCL10eG7WVe6t8VDcHcKTqr/QUe4LzNbK3eBuTFMZ7pVafCgBF8mDl
rXqjpj5M0q4J5jFBBfsSqa8UuSXtqEIQ7tmiJU/8oqn2PiSu/qj+UcAbC/PgudCSPhk6dByj92cn
Uov3b47dlom7EVN1744VxQOJv3lB/12rfhWqZMa/yLkbx/vFIXmjJ46I1eVYQg31diQxGeOlnvXL
QbjryElYuWUEh9l1i/LiyX2QxBkhvnfgXZejIs8xWI2gxTFRIiNfL1VgF83H1+nAGtGPI2noZdRJ
fT/nODqOCxEQn++NJ0h4OlOu4IpcmaNlYio314vJoTxMmaek7MaTCSqs+fzOxvuxPfNrE29DnZI9
ebDJjD9qoTaagclTldv1Y8bjZsdDert8D0VNUZbM2UsHbeOAg0AQNdMvbx64EuKZg9WDAY9azuDw
ew55nWb2UHKAkPgiGzykBV3cVa8cpLP3z59X0U/yB37oU+coh26rOLcGWYmBrHKy9QzM/3iUCm6u
Sw09/upkFIbDjfzNkNab5rmhI4P4pvdEcqUkDrggwpyLWiuh5FEAGc8aO/rW/xtiHni12GR2SDzD
hGgNuOKcowdzGV7f2+o2gPC92P5wvxBHidWYXa1p49DPDaM2bL7AKFLyEmN0/dIXLYYokSHXrpqg
DByPkjGUh8ia/uTsVTdsFbaez4dQ62vqn5+HCjIKj0J96eMeMzs+QjFywbswpRoZITai+DpKtUSu
Pzeug5ES4M0zHBfj3E7QFufNlKV+ovcahOeLymgCkny21d+OJRgMCLEQxFIDHk3WiA9SHTMb54tX
yFLK4IKAzek7p3K9t+uuSVbRWgwnRDY9oc4cV+T0cGr/XU7ri7xqpYai85nvOEXG76SlLdRo90nU
7RrdTKJaPYuCg6SrNOj4kQz1GFJWt+iDI8uOgiLpuFHP4bVQFm2lH98c4C6W0s1ijN/L1/bw+3Oc
Az1g9LofF4LhhiyuoZEB/T5OoQhjGtdB7D+TPgFH1q7hULesP7TLLPgL9sF+3PgPjOYF9aob8Ua1
7SfOOj7wh1nQGjCF/W3N5hBIbyATJJ4JUY9OcoeNt3IotxAeaJ9yaGREus4EOziWSeIABQDI8kyY
lVwYDTwubCDrjHDnbo9SsWPfuaNbWN8wGMYP173esffN6j+U1PAiayP9A8OoWIhLm81Rh5QyD9oK
6Jcpl8NtCglXmX+jSvJC+3g3iaWQFvvMKJrW7c5jP2ulPcMwuvTdCdQo/qPRzP46c/XoOMaix/6H
8X/ijTonMjVrCIiNZbH3JgTZ1WbjrS/18dyFtAtAeKMdXGZaFJly9YIkaoNzg0NABZXFDXeEFGVc
5BmiHRZ2uylOd0T8rQy+ZHRzwdDxG6wRGh8ZuVwNyZb6CHSShvumqCNOESFvWJoAuTEQXbNXnotv
G13lrdcIRtQE2i8ILYpP6cyRsGLSTapKjud0eO7wc5myJWUhq2pCNmoK6SDxxsF7ltXeJHOQ59G5
KW3PhSmdxB3fanxbhjIRM0LgI4maKelda/Oe+d/lRhDpSxbscbVR5Zqgdh07f6Zjl9+y0WJ0zAi2
+fql5d5dUyuWaf5BhZCpZGyZqyqF8qQQRDGd+24xFexxUsC/0/XHo/f6mzWC35jNS0YCTjtDCn2r
fcJeBYqzYLVG92fY2p8jB8Tr/zqScO4LG73kr3V0JtzQJW8JtEBr0FUcsefzBEhc7qdCYECRo/ae
fnjHxNfYAtCl77jIWO+o5AMSuCzdzliz7TrbFeNeb1tcGhzKTIOduIPL5GYz2VvXqanaTR9Xyupu
g4kXsMxL7648h9LuCHBepAlddfSUB2TrHskafQiD6h/LlFejOfX+MxZ13+3qm616mBJn6XFsnI7Y
lLgudqf40kL0d+aAruXbLj5rHLC6gAil/dlwX7zvVIPHWqNP98jAoqg2Nc5K0GRgQoYKBeJi2gTI
PyP6+H3Z21H/nf0G5TxfnTtcUHuFT4dRRh9kRP+GjyzeHd7m/Ma3lUEJju5Lrx8LCptlWoZmgIKc
mBY65zP/tgpVkaKGv2+QLo59cfGXJSj8M9pKx0+Cb3fN7xE5JJN+WfGbRQoTvhs7BVID0HvfS9BX
BcJtdEy/TWvpT8/yIfNZscILVTu1Q4gQeuruQDvhalvx+M2tNpmAOs6jXjSNTq9eUFJkTTcFxrZL
rSSp+IDChohDjqiTVcr5xj/NLU8lWECkqe70ufJG3ARwcyS5214zmnRUIomYCGl2bbQUxq6PB1nx
KHfAEs29UogUDPcc8+RP1b/nheDFcTwigR+zW7qz9YD2Oj3HNoVtILNLSBqwA92yVf3/5P8GVdi3
DPJ14VHnzOEiTtRyGXlZb3M5Z8iWNn3vqPDLAf1uuJltxNfmmlj/dhv2cwo5PKiEXVJBOO2qgC4X
pqwjFcxXnD8ACs92IDHQnWaRmlnL58T3ycxGEmZiHorZXj6s8KedU6BcE83hdAqfNGQySuzcdmzs
SY+5k2CgQ//8/y2EQaF6ErkIIQYyewcGSr37EZttRTrfru9G+CozmQEx81THKvyHgmzToTzZ5LTb
trcXBYO+smYhY58Gn/zwdaXNWvdy9dZtXVM3j+vTuKdmhNxZToqW9AIkEnuK+NBnix7WV2cbzHg6
yoou+wCrRDEmq5nr7DhMeylupbP91wShudlz/XoBuIVutJJctc7I8nJavbwD49qW8xIp3AcmE6QA
wDOU3H/ecnNX//vnGNjjDKqDBTGC+NQ40uvj2HGXv1k77U5IslK7hhzcStiPvJkaKThGutjhyWNP
q2z61p+hC3aQ52OttLz3bNuTJhgSnb1bGLfZPF/mEqsmEo7VQwjQH404Hf9xZZS+DvNEZU4jSwm9
MQ81PjLDa6dsfjYLczCd5tn2gRcjLHfMTqcj3sZZRvwL2Joj+ahnHEZUcD3WGSbm6wmI5Z5XriUw
f+wJdlnSnnLOT4FDmZ52ZKvhjObNpauEHaJ+4hqxtihfmNlrySkBNR9MidqIMkJ9LNcmbRjYk+cS
E7i4scqZ1hIx/9aYT8pgwSDW5knAB5dkKJXYXkPxTE+cKddb1IDOfwAaOwYWvHLZiSBen3Ai4/Ti
2gbS/TJeI/bgBJZW/180C7kUWuylazjBXkOf5uVcsBL9hhyklkPXp1tB5ZURDsmysbN5dauNOTmp
ooeglzBz+hv+Ccu10yfXVntpYhgfD+/6A2X2436a1fcgs+qxK0a5E+gieV6QAZKsMDeXEtDp9LvP
pytWscw5qLajvmNHieylhrI8/lTlkOXVLIfFaG9bfRpbZFOyywogiEBnUON3tBoQkdlGaywyewao
TPJAqur5ZtA6etI6RD+rooYdYA473W5041+cEuN5p/WcGjv3Af/jsECtWImeRO8msOEou6Bkdjcf
F9WC99kbb9GBYc2ycgrecgx8cI1xyVUDmRD91ZX6PymF4lgLk1TZyPolUK3vhOi/EbQpAsPo6lBN
d3RX7Iz41ToejGpvQjkQTCphmGlOJFEA2q89IPElY9Th1Dm+tIvRupuYl2ec1y26fPcQvZLQA7ss
SKIMRbSa84/QSYlHjmCoZC83zZJQwZaY4FBt/2LqQ0OwwH2Pv4OPjEpkZt1oPyHeKNz612COtzgz
dN7JSPn5ukF3vY8zNUs064ZpXrjsHiqQH8kPnuX1fMaSsQRxGfB7ql2at7+4hOC542CZIcHCduvs
4FPcJcX5xTyg0tG5tp015iGLK5eLY1RGdVd/eTi6tuomOWKNnOOIGI/nmKwLDLXKv1fH18CZsg8g
Xmp2UVXCOEsjSKphCbx7ZUr+nE9TI43K+/rt7lADufwMYVLpucWejVJon2zqbXq45iUjIzFybXZr
W1OHdIUMh8oUOnzreohsqDqQpJFOelLxCP3QLC6yrE6i5rL3q9DNaf4147ug2j1Wl2PipndE3ae6
kBwEjFuU4II9nSHQYz45ta9zNMH1C06OQuCZivLvFBUe6QDG45VBPQVq4KCYv5Or4agI63coIdP5
dDDFmQ2lLbOTSpzEsMIyCqF+gmctq00ja4NJrPyLtv5Z3B+aU7UYf2nT3/K8Zm45DawkZJ3Mr+Zy
WeitVWOgLPCFaJqwkWlHJFkULVEDjMXhIFyUHRmf8QHLnDCNNDqFg4MalrXq11bDZfoyHT59rXrH
o4vBGGp2M4fZIJQ21rRGyQoZrUm3e37H5cguFd4v/WvKhatgyg2e60ylSJDQ5NOwaFSCyxi7LskV
WI+GbDNhLcGCppoDKCKKQwUVQuzGTuQ8wqguPx/KbkcGlI8AvSrEvAdwDFHWw1NLUedRUc5CB4iO
BmwLpLlBs5SPxYQpUVx325cYJkJHwz3r26birOFc6lFIgP12j48d/bKY4diG9LPQlUh9cVeoQCrT
Y4i6ccIMUxU2Uc/2kqDzqKaTRjxjLmQkwfgcZUfUX4BsVl/09caA35ORWpsRzSbXenJvI8WfdDPW
V4CcH2gdaSJR3eOU6tZUGnSGuwdggyd8SRS6WoQvihkogL1zSocNavrvuO3WVSYhEamRMDypuKYw
4u2Zw02CQxfwiDUBJKR6ya9b39gpVEKBuALRnaelv7uvybmguPsTR76gQr1QDjmKGSgG7dAQy3/O
W3vbmpn0yAAfOJ5fzXswglMHwUfqmgy5KoWzjaYw8m64BxVmCMe58+ni9QgyJ/ORdelNCy75GwxK
MWKq/Janyyhjae/wdyFh0sPJl/Ls6oqA9f849e5VFAhkVitnV9+hfKM4oprsYQxdqBuUJAv29jtc
o4Ar6p5bKWfxOem4LVh9rgM4PHd7W5mFmnVxmCFx6+gajrwDI/VHcZkAF5kiKMGNRggyrY8ZuR9t
uQULVHdnkdQHtI3BG2mjDk6f+puLu7ImWz4dEfWXIuu1TA27eb5TuGYQeNIr2RPLz93vgdY/wuFM
oFe+Qvm8GC6GRbxbL2aY8RuZISLpmtA+xRCysBgTf4yd9FSWQ9ajM1Kl6gE60n0CVi7CrsQp127q
apHZ3R5UkWzVp6ZDkC9e6DCPf4sGZqhJ9S0wFg0MpKFPXlqWwJACT1e2AcJLuT/LuhnCt+MLMjgB
O/ElJjKqpspIpUp1sLMyyoI8jCCZEMzPMoC8FjdxeeHjb53i/OTucZ2O8eywjEH+1A2qlF/cVryN
olmyS3EiSVuHnithIDKt0UbaKbCAadS0bDSwGbKGLdG/T3/4/Gr29vsls9Or4E9WNzR9SJh2/WWV
v2E6CtMebEAvTZNBmaQpT0kEjxaCy808g2VH3+hnlU5JRiRV79VsA5NK/zsRsWGEvCOFCv3kapWN
+DANsDDYbaFG/Wrc2Ha6LF8622D3t7S/lzgYaezveKV1i/rVrBPkRyE7lcjS2lmbKpP1Xa5kfysK
d+HPylGPeifYnixAtIbvtPOqz+Vfr8sb7ai/hrPVT9m5gn5ajJ8CKV1LSKQ4tBjI1QhjmBugz678
Ha1vxcypJQwZR3zVIjimmYvfyX3DSyk2YVUvoAX0+1yDZQTAYqsj9MDOwClXV6hmQIcuCcF6SYl1
yLhrUDgsrLLG3DJZh5Nbdu9XttRKAQ5oVQ0QzX4ZsKPigpiRHhPfgZElT7Pl2WLWYiT9AWg8ns7P
2fxsfgvQivNErkfezuzNpoDUBhRGWNY0CIxd7T+n6AOnxkF8mpRo4BPNFiS9GdO4NEaH8eB2hR8l
E8ik6H5UNQD02jMrShlToBfb0Xi9fKaQi78TMUGiOJVrby/LTLa7egGMl9w3ANKszfdY21bQLltV
3Wx5Ni3UC8IcfAiY4diXjN2rjDyXWAW/n0RQcF/s0Uo8N6BJQlzBZp/W0asN2IG44DHzlUpBkzcY
pOG4jGSG+jRg8ucxYO/CJqsun6KX3h7aitl36u/wRJDs2AnmN2XCeHH+1cCdFnFYqD8psPpmybV1
q2+Yyv7vgVwtOdkUvMvXR7FtsAMADxup3035zK3Tj9LwTO+Jjx8dQWdR2Ooyw+HZOFocdawQvkkR
QRCQTizawHOVGvNblHLBMZ7NwBgH0DvPeRhmt1G7yPwZx0JYmv1YB0R5boyPe5Qxz1Y8bdaQPOYq
l2Ro+i0qL6NFE65oGgJuJ9O/FqyrQFuy1ipdMoxf3USfXhgsm806f5fWDZE6tgaX+8BxIjTogt//
h/diC7sRcnFhdl0Cz2EqXas8wD/I7bOFNnIlYq4Ux6nNZCRhWrtShLexotL+4zXXfeEw2O8th0dQ
GhjacmpZDqk7BgXR4UY9cOzOWeYJ/n6wYh1M1veFo9AYpIxFkusaAEEQl9qssfmfGWYtuLTe0fhq
K0+mbWIuqTbL5DQnpdqj1rMKeUX33Yk9hrczo70gWeBkXMq8zampEPNEaBooLRgrGTuwabVW4hgB
4QsOKiHeWkbVow1bguXi6HsmwCE+BD7J6aMvRhKx9pLZYCbvrFDp6JCzAkq53yA0VO1zDn8G435i
lbtLReCmGDbnIwEXJKpN+q8Cx4/5cwHmE27O0vf7yeU+s4WpynQ13A9DkTY10vliNkBFg+NHGOoU
G8pBXvVqNz5Ewyj9bk4Vt7xGef6Yt5muAiV78Xw8bXVOA+WElZ6zUaK4fMVocvoSp7bLRDzPlJoW
NGxQIKU/4nrqGGggeIyTz0Z/MzfOZm8hBFue9XS1OirPTDq/o5EhAoPYqachfdxzMoZ0XG1+V+3T
BL9xiFefKaBqmMb7y8nBCtcrnO9J2xWVI17FhcxxXpXibajJvKJq934goW15TT7XpNzXGp8ezY+R
kGqQXzY8QUQizkco5iK3YNSpGJphpkHo9vRELcG4eejlYNn1L7s7WSvIn3FGFKdMUEh0fkios6x1
1dmFyD6t95ANtncoMbDC2hhHXmpToCTw4Po/XtlA1VKH3cLlvI94HaMtgZ0gLTZWSJwgGjkG6J8e
5biItAN8RkQ+ZOSaJN2rhaUrKyxMXdjPjZldldYLRQkxXXcm+wfywnyBEDkwl9Db0ZlDGL5t/42m
FT3Hu1de6zkGMmLG2QKW13YQVZOmkQRrnjVi3q8MmEwm1VzxqVHSYtm87PeZ2X2FyRsnA928ldvs
m8QhaitCSz9X2q+cuiXgkVlcs+XsbFLRZqTc7CMRC9F6Ge1rLqLYeFpa4jZEvoCTkGlW6mqGSNhf
OfblMPWlNPSFIJhd/Ia9MIFb89J47YOZjWUKPB0WbndogVde4oUbas00YFGBWUfyohgxmroJhDtQ
vPgMRxkl/eCYBrQQj65JKJqH84CRsB86RCxEhevJBrR7SlsV9Ys4kFiSOtnjVIImPSJkouaR9AhQ
dWyGCtztVrPut55ceP0EF3n2K/X/3EtwJXabVw281wF3+6Tcs4E9Bs/nhuzJISVH4TX/p85WUBkF
+BM2WOfF3bEcfFm3ZRxl60fQssEaKVfu+qRTIJFzlsDnLpNpoA62Dukt+VQhADkdLRDG99XuFuH0
SpLRFOgO39BCeY0rblgha3oaqtW/eeBrtNi7Ag4Kq5RLKNd9P83kdklmGbgTzjOG1ypuWDPqHId3
d29ra3FRMlOU6eJ8rdB3VOM30iPfPN2bFCgowFyCD4pUtYCnUBp9H6ZMwiN+8Rp1iOrnllOl7Vb4
k3uNfekk7706beTYZWQNsRqbop8Lrdpv+30X4Gu/26+lHAyNDmad6A9DPpFeSRpnVnVM+Yhr8VN0
VafSkOX1wTMp3s9OSj5VqqphrzkDpxvgRavJtTgJLLzCDx5c2ckSqYp079+BzZSv89ikGxklXKln
qdd0nJt2yJdW5SRWTewO7+y4Vuw1FM8N6s9RYwApDVaGtQwTWueEKsP37puDAtQSufTcR0kr61T3
su1/Oc9XfidzY6CnuuXMAuIM3cRUMxPsK/pGTrCGej3/xQCCKefqK0YdF6IYvbqXktqpHFyiCXsL
0qQb0mNkCARBgsg3AxplXpsP7BkSNMenJojof+liz5Ajm6CbAaSETZ6RcQwTbvUb65AOSHVy5vNA
2kuzDz2tSIwjQ5oe+inhIMJMycBH5F10UWUU6zInERKuEvgI+mXIYtc89S6iNAYlY90kawwF+5wp
TOe3/6kofjfqS7lXib9D2YeTIRRxfzOVxMj7VjVViCU6vHBLSFABtcy5WCK7TiZZgOY/o/1N+s8t
UIWVVVWtFtNYwGj37K9Yp1faz0BSNoU9hvzsJaknw1lR6KU951KU0WeU2PiVInRmOzuVrY4QZW2b
1Q0efsrOMykhMPbNBMvBVBj3DdnZYLqv5Wub72wFE2gAkhiBYO24rPfXjAHjGrs1mjS8GLDTqEmV
oSfpPkM1O0jfINylT5xIKtYnc73RnOz6u13nJVFSntEK4F93Rka8odTto6C9si5pdz6qHSfCu+w3
IwTLVp9gff1USz50+5Vf5uAj4vJnz7aRtgibAZrfPaSf0OqQeiJbrRX44cbf97zQDGZ4XvaMJtzd
TYzAKysIR4TW9tBRU9jizomdErNYZQ2a9l5+eI/ABHZIMaTgkkdB9eco3W+xCuoti2O01w2OuV4u
st0c1JBiSgkLjg7tnwEZmjfkKLO9SsJUuShBhG+304P5P6dY/CIKcMA33szEdPo52ogPdosPbDtu
LeB+0gPs6r3Sj7++WC5r7EO7zcZi6NIMuRu126FRqXpn6HRGp2YE4+rm5FRxLMRAiTDm15ilY/4d
GQQaYJFdNdWfI7DEo5D0RlrqIBXRaJ7c5uFKA+CxFzq5A8RZ7TmIKhrzMGl6iWQhGjv+3sAKQB++
Ag7CwXqPxzPhdJITeL03q0L0dmqEgTBtJH7AsnvcV9isyvfCHw4QnfXe9zTwCt48o6tt12TjDq67
k9Tuiix6A9kZMkjzmPq4rkt69f94rN/Lm3QmIVrG40KwTi+yutZJ9IKmYz4EKz+bcdfzWmY06mwO
i522U44EF2w/F71aDkmYAfT7cvHm7Nm99imHSii08fJAjqybe9B+Q2DFgbGO8Y6RQVV0lJHNQ0B3
fkwzFTkKBfwBpWOb6wF7C3IX7YL6VvLw5Ik0iDqUPFC1cJWqfBpW5vk+91e8/9QtOWzVMsy89v57
56eKKEHoP2gmqTf1LLBNkcS9Soqq08SC/YQFOJ4rqdITTRy5VVZLZzqYfR1tYBgxrYk3lXXNCJDj
wAzBTKQI+rTfkfyhy3+x7wnzawbB5l34fdM7TeTAN/wvLJvq59djvTW6xxFsDeEHeLr6Y0QNb0RC
l5VBVCBseVOK2ckMcDn89wKH12tcj7E2Q26F/Twx4ld4Q8U6H+Y2T2nJ3UVsFVTY7VTDJiEufoWT
MscNWmG/gntCqGmA+ZO5BSyZtPZm3OV9iFQzmEi/sTljDQ3y0zMMMzmiZ0X4GTAJIAsQD+k4bhUF
eqPOG+j0EpLwWGZLRZoy/dA0vGFAwv2PD9WrK0YkrNoMQY/+93PEj3VwK9CB7g0Dkdm49Diaom+E
Du9W9bGgESbRkYfGgHCDu2F2CjIdk92/JYkEOrYLGtLNDQE3DuCWtDUdXzN81MxlAMh6zoXEKSuh
N/fNtyD+YTI4tsetigXn0uV7t9nv9TaZ4y8ZkLoT+ICNYgykhiR0jRP8yIgNRWZ/9I1UwlWQ9MCt
qJAficrmYSdvNrNJ67jbLqhDZHkiydIonMiZ4gbG3quNAb9nYlHnMrN8F5KVLH+BbwEB/4pm2WIj
8Y17m2n32+yBPpV6bnjAYzX+D8k4pX3CL5bG+3o0NYatxJPFDg3aSxyXq9V2tj6H6PgxXpMSzK4x
4R1of8iPcUXWUv6QPXJQmIqApW+Gvzfd0jkt25SKdJOGYqTOKda3NCctp9ScNpMZJHNhroJZaiuq
PKYTqyOLDAHMGM4a3OuNnZli0giIqllZRtHNoKJod7XgcKBaHCTy2Qdsm9wm0iXg41XGz4MPIMrd
cbngBqlYodt2YTwxQtmvgsUUjbxDpB5VTaopP28S9cqjjlKbmnXdz9LgiUs8nw2kHWlcXrYrFhuU
+8yUkrRWMb3sf9xYbC/yIgvyLBLQ0soWss4k8VYCbuk4zJih5RC4qez905IfbPe4XILJOcD9LNMF
u1qj947FJ4ABoOF9ZfNP97EerE0jCxtqP1n7HZTT0H6JEbWVYuUWUE6vEHsyhlblTL2wbnMyRnml
/zIY48/0qmTJOubPY8+HYHnhAk8hMhESw3gxvMNSUDis5N9CEDGpKz7x9jSwI2GnVxMTB0YaTd5A
eWRraeO06WX1p9OvC5geXLqgF0eAE1Ld85Ix+J46j5eFr0upb9H0/SAVVl4K+u+LSd0UCka8pu9v
P90wxw71G9y9+3/69Jbd37AgiZ0dRH2a6GD4enepY15whhvB87yePAsZgQsq9hw/4OOS7UmehDPC
9dyj7frPhjBoanIkEVTNEv56/ygtG3RKi8YjT/AquInrR14zNGe1vYgqh4SdUHo6v/ZsJKAG9Xs1
MdMOETzmcn+2mgA34zBKN4Z7yQ4pjIC9bIHSUbDANFW5hEWhvE7TynLkU+l1tJI7VW/3mNeovO2p
D0/1IS0rGQntCcG5Yug8acKpBennvthc8z4D8Y3eNQhgDILANgvCFIEV7vnauR0Yw4u0z4d85STC
pngkXpRPWv38XurFE0oioHO6M2sK+2HV+/5LSm8gEbr9+KFkgq4ETH5q2GHLdyD8EzF4kS4ows4U
oa5pd8TiQ9Wfs9L55ydtLkO8eKKQA+5WEEJ3QgacLeFAcl36Lo95dVbXTtY39LnPNssmYRbThtH/
4gm1vExhyJw/SAFjTvVacG2kPU/7zG+4DSvZbJ1TuxBF3txMxFLaIAsaVx/UsIpT3BHCU4bviOC3
oUBCu9YZFJ68zGehv52DxxNhpNccc4ts9xdTsmGZb2yL0TMfPt7fnDJJDBz3JcK+tCKlq5I8sxBY
Eiemanr9S5ZJhzf25LH4HMr+ngNQDtLsz8XY9ho7Jiue2FkVlfLgtkY9Lt0kR2WLG/KHnHpf0/wW
uWVOoyfG00cTRh8EpjSIJlh6zhc9iUHbpwb4r1HMBw4c8ucAJDhTvIR0hhdBDUsWQsf13d4IuL+p
IFve4LtrBQ8+wtl5LAYhrpfnfrzIK/LZvhKjmPJOD6urAzbSUIfhqjSifD733XEcKXhrHyCm11fi
hgRYWql9r56EhKl3jgCbCYzXwpydGZ6ZJa0ndtNXVJVodSu0foBTK/gL2+dx9yKeNYkD5yLvNAMZ
5cDLL5BU56upK/rw+8I/SXKDaDLOzafvzoVlaIa7ciacs67+VKoNcygP7J1adM1v/g0/Yl6rWMdD
2ufq7RvRXw//5NiIqKond9K7dW6BUULy/ORwyjO5rjcWV+5f9Q8E0Q0haZGcVU66aRYXM5kewSVk
0QlJ/tzQ8Pb0/i2pirKlrbPmpC9PgIKPZ55Xqr2sMWMBQJM5+2nqlPh0eh3qdrtYa5WzE57ETdbK
ae7n+VSeqKeT3MiU9p8Y+wx+GW5SamrH//yosRQZMm5snt1dKaphS7HwXns3I4zvc4trSKcaYpLO
EZju7aa7fjv5tqKipcuvVQkS5JcFtDaAjK5fNB4Symg9QamXjiENKq/KcyIvJlxBj5206Uur7C9H
gfXwYwws7RJbvFZX7wXrltWKLjo2wg9qOYIGxTtSclpnvUfoOV+jDLMfqj1KFUg2s0s/QdmbTNgH
4UbOeureT+pcbXS8JfeW45YPHr5J8Dpt8+rszZKONCJLeYKLNrmgSCxCBYAFZZCs0XpTDhnoFtqn
YtlI7gsHKwT3fvlrVgct7cm+gDrrWX9HavGZ8tnGhTyQ4LDpykMidQSD5KtFrjO9NAd9p8BgoOIE
ayHMOxmtjI8DylgzfOjZMM11G9vlCsckqPrl9vxnnFol8G0DFWnbAcewp40PE7SIyi0Nxq/FA6uH
/2SHlKpMXfklnYgRIk19W0U+6wATPxuUvx23+ytqD+ZP8U+mCBT4VCwi9sdnktGjNO7dSwfSLGFa
HvAQZydm4jmuSo05CWUEFckpoE4yH926RXM+Sfm9XFUtRbY9DkJAq2UZ1T5aTkVgO7YcqSV+j+xz
qzzIr3Mai5vNI1pbP2gCgjFHEXCUu83vzAWmxXkgycVYtndShE8zjQo0PwhQsriXsQs+lzkRbT3D
+Z4PuQO/8mba0hg8q23eBPUs+lr6UIZ3VloZrydk/uESCsdd0wc9S9YxvhMz+9d+tHqfUymiDX9u
JeqkbaPTXPlH+aA/cCTsDO3IJnbJ60UnNI10oUV15VIKkG0D+GX3pAtcz4G5GLFN6gMoUxF8WUSD
VIKCzy9rISAKKDtjc4Yd55BDzCE3ZNSFkHTabUMXaiA9CO6Fk63hu+kzDhiHq2hUkPxEJoxVJd5j
Rp1nFUwSW9m7XlBabqsi0H/tAfOmrICh4XPajL7MCmwbeYxc2g7txnlRheY6L/BqsqmVZtcz4yqN
UyRMmGwGD/0ZglYLt6qGNo5OqE4yhMlJ3ZTAo3H+bY/LKxa2IIeukIyFNLKvCwEVPYPet7okXJn7
ELU3YqKowd5P9H1ny3+M4/lc/y07XaMbyelVdACQDzsFhtRTqSFnqL041nMAXMtHgB6EdTmx4BVU
lGPGW5D5NzWyQp9LIonhn+Zkd2BmRUhwAiTNkGGTBzwhNj3p9PjRGEHroD6RWs5bLkZpF9Fzlz7w
77hJcdMgMuGZQK6TjUVVUGQbeMds/ph10PObiF/gj/v2Qly87TfQ4bpNdoj0vRYojSbMsePwUWqN
E0716SvwcWtpplJQwhX7h2TwH5+QxRgvmH1rnmJbHCf6robeABQgy+1TPUCcu/B6firMxfkFGFA7
D/7RB5cfTwEniqVIizrb+3Ys+Epxq5fhV2W/XMGOwjCd+596SirX6azS/maNLmzIhbhjNpzJU3xc
EBU23hWi9X74DQv1PD044hUjM3ATx30t9ppuAaqfhBse6pdDGXqeGKz99ZlwgDysEtxZUIXYm62a
5z5f82jaVOiOE0eatoZlbS/pzKTN/KkUJO3tyUc52yMdoP8xtVeTVhsdyqqz0sRISc+ZVjxGOD3t
OmCteXqXp2SSaELi8A8GtL7Sq51Xaz6/XKB1n0PUJdjQ3XZDLciqhdZ2n1bqI7plyylUlgVjcMWT
lJ6nshvzfy5R8of7xaf4V7bf5aM503QvUETgsv/AnFpJPc7Uzf1hGTX1yk7pHgnvFWEcs8EdkdYm
dLumyaKkYehWEDu8nSNHBFHYOpGYHjsxCDZyK0piccJD0i6kKKyV6ACLv3XqlP5D/X5vqg/Xy6aE
IdLECEexSgKpPb85GBKUcYVsV7g8bfuOrITx79x7asxasuFGAydxJKmxkAn0WWRvaGywjT9nUPIT
Ap7vm2jXBo3grGwvLSDWreVyAsNZPHmqnd6fpWN8HGsYFp8eu/LNLCA9qU93rwHWGiOQikE8HZqE
ax3PzwxX5CfTyq7iaUpL9kilMSj/5YLS/6NO8XRNVcQdPV6AwLmf9yhD3gjNrkXSEm7kkG7YBTwI
aDZmCqFM55TtO/VoLLHlZWj412eX854YLFJVMsa+YZkg5FAhZpDICwvIUm9PB6n1UAdSBZFLGfc1
qFlBe1LuQL+XNpA2ezyKRoJ/NgDLDUdX6UFzgk8ROCuHCxq8JRoLvQb44FeCRznDkdlK5BrLWCKR
SD9KALPB4+XimZn+swlzYzpEGjAnpbBqorMhlmUyoyTTPyCtgsVcafpeR/uwy3workspyCUb3x+0
BrvCP7+PYQbkSh20AHwcSuPmiOzV69zzBbFJWzZp8+aT3pr8wRtxh2gmrxEeTi7eL/sPpw5Hn74M
+n4UxOrtufyR/ZcnGu0uiarim76cfcmiJ9rns3Wn+Ygx6fI3jybGFyscln7zfYwt9BWJoGT+CSkj
C+0WbJ2QKFSmfGVH161syuhiPLzB6anoictZ3jqNyrXZzmvMLusnViFmPtM3K1OR+ED2BcVvqpV3
wRmwBxV2TOFecfkSjZEgzBiDlcBmnGwvOYFV+YNJMGqT1LFuBzCUKmCYsF4eMk1DuT8pueyQXGDi
iNcz5/aX8et0cWX3k09U1eYA/4oSYJVWfXghEgaUqeTyyymPNcp8X3rv+Vzm+M7pMnNy8MMd0EqN
L6jgFij7MrRuC7vpZ/SthhKyRpMKijLxyRxZ9/NkiAYK0rtvdtjMXbxr3sZXnaQ75UYZTt9whAch
nZYT+AnFktyVYcBWREGfBFTzPbPg0rdGcOGEEOdJaRhrymRUmyL8GTwcnCho31feJtLcLQKFBVua
nyv/Ql+66Nw0dFiNAUv3RWJ7go05DYQSnjbUHO0w95FEp44qrEnVmn3M2k1YM2kSC0XfsLW9VLLn
XtSPyFILxWujQwaQD7g4oUc37OZaOMKUNgcvOIxi/Sp2WjV42tSvdZaGqshKYAMZsIy/LHw49Zqd
k7m8oV+V0W3o7SP764Rf3NRvJDbeuJx5/tcufcSBc3z10ZpnJSB0rBvTFgQnEqlPSE1EbBf5i2Qx
jkvkr5QAoTUNKgHgc3Pxdx0WZYUOm+M/YOu6y8FB9nhcDbZDz1Bi3SP81ByXuffO0NriFu5FKW0R
nZq7D+/W94+0j5A/5v97zM3r3VLYK8uiw6FgltAnPyeEyPV8IEiAjlYP2WVg5ZxlmTUO0bQrOEN+
ni3rzVyZC3ib7WDiKOsQbKOFvqaWbasFXXkyFUdxzk5uoLoJ2sRQI3sj/n5u7atMctZz+rrtmSxB
ZHOufTmt2jsYyjKG4ZOgvRPLlbpHwYZkn90U5E8/Bgbr6kM3a7F7Nn99D66KYRO1gbcpyO73dfbh
h/4wfcchAIqtoTcxcMbPmVKe8FFh11wTsrIbSgbgbIiv0WEHVO38ym0ByS+UyqO42GeBj0Uz3gqj
JOY3+V63OjndjPH274cYgd7hX8od/eMqnLyFoVW+et7MoWCi4c7pLxFUbZd9BzBNurwN0uX7yZg3
n+4xMPQAEqxOW4xVRWwKFNsHnACMOOlOZuGCzJmQNq7vRg8nhcXHh8JSWUEfXs7q8+2ztfSnLuGc
bjSSm17/Vi4XCXQ+mmdR+1lrDZP2qA/CCH1aKyNnqObn7lH9z913vJ34IGqQozDnrYuCyW4pQvK6
tl8OlXteIHn+4DBsb5U2KlPHbIsWLFpKsOjCDkiNYY/cAJW9DV8ahMJ0oAM4wcxycAQQGlAsUdyH
SHpAmzXbrDCqjwtTUXHrwibsgRQhqJa0fLh9muBj+mHU3sOQse08ea2oZCm9O369omE4rsg/EX6s
zhrfjBGL+GCeV4xvL2zWQOluvbjp3lhq22NcHPLsrr9xxAkrzHgeyDm+Sw0nPgT01hZVQjgsNozG
VH6wbEpT+Bu4UHASjZjMgCzWneVp79Ac+Vpdpu6iWpEp24/S9MmBm4dvsT8jdhlj+lKVARKNf990
/Y944e1uDjTRkc3LOg4m9mk2FS2kv3fHfagdV+YNw9bN6xkerzkL2ek2hX5Gz2L/IjepeLsGzrI5
kga39dGAqSrbl/BfgSRH9Qe5a88PdTpk8bEDelfDaPL2plxS0DEnhCx0jyf6I404UNNhAyadHEyh
7wWhOsAddNATBqg7piTpPkOLSpxHJXyUEq5eDIp7/Vw2tY8zPTCsW/Q+2tiwvJBHHJitvYqkX5KS
Xgs4fK2kQsszTW3+oiZM/Hho0pEzixaAVu/0u6gIjkgPi7E19KiPiD9Qehi3SaN5sb6TGO5P87JL
mp3KJN7kCwrMPpOkEIZ8/PQzTIugwYkF56gepgkN3mejlksRlTQC7Ez/2W28dzRLqI9Gz63xfT7a
Dp62Lp16y8rDjvSoCgnfdruFBHHFcWj7/sdiOqcBxXNQxQOZkVDxsFxW15VEDKfGYOZRGWXx4vym
NsdnZKmU19PoO8FVkyoMd+HtSbbhnD7+w8cn7QBjLcNMEHdYsQzvKJGfFxHCYp/tkuNX8E5C75xa
0x6iT9k+4sEXnyUK7sKVCX7Y75laBbCC/v9KYsmZvysvNA0kl1XkyTc/puaZnxiViELa0Zvw0pkc
aukEdngZUA4M8Ez0j7JcdP/rpZNpvYIono3ZeP+8ySqHQMhzLgBPbLxIoYlO8yK2Hz/AZXvcJT7F
zeIsx2TIBQV0q4vgzSmJo6sNaehHDjDZLFmhjeWPqfx3eFcIRYS6X3Ck5ya0+B48vyw/5dJtwXrR
9UKKcRtiFuNadhBB5QZLlzkH1eJvZTeD5JdkpvHSOxiHsGR3SUOzWw2Vekynw+7GXZ/0qpU9VlkS
Ii35F5tQQlaw5gJyBkN23JQifYTzoh/8qe/rudtkqwM1LqKg/qCkhx51D4i61r8TgkOoE2u8S6A+
994os/TNPeE1tAgCfncieiK3vsdzD3x0zm/XUMPVU+FH+eU+SAGehFwUwcTmNMuN6mEdTFMzHCAP
ndCvik9wrvoQuCQH5HTfW6GJ3qJdzgD7egJU8G9X5QQdfLxhiLqAMnYYXy7aMxNiTMU+C1Kvb+vU
XqUpCNuLhHKpSjG98Nr41NfYQfJUPvbKfbZ6KSvDpKDI+7VQuH3G+ejlIVzKKpCexo/kMXYitmD8
QLL6IiW5vRBZNPAGmuYaxDd4ppwGBcPb7QMS1hlBLihd5fM4ZOF0nBXsIbR5i/3xuAhyFYruYJ5Z
zAZW3KPUcmlEe3Oe9ubsj3/zjk51wHNrappoFKt9DTV9XNajw0++ObV6yGlxliS4RyoHU2XOqzk/
SyqaqLFjloM2VN6xwy8BPL6XomauSPKuzIDcVAshwf8DXiSsP8Yi/iAApXR6ILvHXwYGRrgRH6vB
NIzZvJPWNaa4V6WHnJmu1jwGrnBXbc0GifMufCzv1k430w4XZxGQuggOXOPkkRp263RI+SgDl2aN
NYOmRat86hlJNk9QHt/+J0Qxilz7PDbkPVZLilx+vwnH+uvedGXnmnmG5zJMHAWa2PVODMUOlQ3E
tjALzq/yN14FYM+bXNxMT7Fh3F+LFCRLIGJyxnUfXY2jDLm28P+2DmaIvOj1s99G4LooCStc4K4z
0lPRxE2n0xrppoFbAY8Nz+mzqko7zy7tqPQncGqYc+/O97SLCfMMfIhrcuSv29r4rTda08AL+a/7
gCCLmPKfgGgc09kV4niQ7HM21Tiw5FMSKUYyC4e0Bs5CFsw8lqKdGtOw9EdakwQ601sveGkl6Zo3
hv1z+L1+4c/fWgR1VcB5kvJWMGVFDxIYu81hC/I7ePq9aDSSW/h9l/vgGUZj7CijPHYbHaEoy8GU
ww0SaOi16VZYltTP/yFUyccmVMEw56jXg8viCepntZON0depb04S+ty401+JRh10XHv5gmcrK50Q
gm8I4l+FxcywWH/nzBqWcJzUQUwOZ1k0Gfd5TWe0CKx5KRuC+rhND0u5Q2b4Nx59rsyfANK8Djiw
9LhzWynv6FziOa50GA29PxHPGBM8UTRBtIrOEHbGpoQB0G5wuc5Pt8ub1Fx2hJgGj7+kRkZsTOQe
HRn/sI4F3MRS1FUvQkI9FhMC4BxeUfJut5mGnBf7uia+JM0FHPYZxL1D3MAFQp4G2FbEbXb9RzLt
1heMRPRzw6zsymP9nukyfFx1D/l3etehXXRsYhfk7nx75ajT6TPGF0IpuZxAJfub7RyWLGyT0aIX
3ZUp80Ii+DUpbqK/rHm9EECvLaRmx32QpQelbpxBr5bMEy1r1HW9OhvfOG3UX+DKPWsZEPxtKqGB
T8dLArh8Tt24IXNMjZaUiHBhgKpCGXWrctWm5VG8Oxsi9bVVQ6wjplfjaPk/044YgPjZcoG4b/jC
foZy1lK8Y9h8fKEMrVuErmmdhNiX7NE02WANWv9vDh+je24KIBxY1T6Cuu4gwh/kXDl5bHwwTv8L
YP5YFWzN6clyl1/wx0JCeZ1LQOnq7wgITSCjp68PrqpG3LRUgCAXU9TWf2dZ24BSX9NX6gu2mgkq
zVi15vrrlIiAIdYG/VO+6hWBgJYs5GlQeTK47B7JK3e7IwkO67PgUiK7Hdzb1d7bKKxsYJc7JV/d
LLOQ28lHcFIS5E8TSVYa+52wxYXSfiDjeBZL7ZWDyYVut446yNFHdsYElsdbknGdUz8bFAYw5Fw/
U6/S5woKDok/AxJRGNjE3hzJgcIBOXAVnungrKh+NObcbtTlMGTKP83T4NcVLJK30Pee/otjOWId
nI5BpfJjJj87zdsM4YU8DqiKMFc9rY/vx2pIWZc678bpbCWmLYDj0xOxour/bX21UiSvoNkW2kJi
J8H1osN5+oA8zNqanA0GuPJ4laKsehJOBjedvJqyf3PID6NQ7ltajhs1NJ51tIGksDKFHVZWxAPh
8uYa1In2ktN5ZqKS/PweZVUZdwo4R1MmrVqZnGgHVQNBHSLpFkbKxLh3eIxQ9SJhcBf8UFVTGQ6H
W94JbgrrAJcibNcRniLzgqmJRQqxsU/DPhRBk6GYUQcFhS6vRODXxMDuSlP94hTB/7sPYD+b/TX3
kfSwfSSCLNek0rzcC8Ixza904byvfih4bHsv9/6xc1cxW2Q6fDiNs7Qza5cZG9FIJxOVNZzNNF7J
il6lM21TbfHX9dVOjRQpxHt9BLYLT7BO4FFpp9M52SygtLJIUvVpEbqv/Y1OguGa5nP6MpZXSKPW
JAeiquwALjFvVYjfQ4LkcInHyBjc2vMIGE2EChHgw6CatnJHxUxidG0an+QY+JxeHPvjiT/8WbzL
C7WNbhBzmGlVGpdmhX7HyPxeAJv1VWYWr80tLmMxXzHTPAorylsjjddOmayMH9rLDB77j89XBKsG
UakduGjCyDH1/MOohv1YRJyOfY4t8KVn02z4dPqql3ATW96jkaubVr0SQ5tvLJe+I4JwPGM+kiIu
1pJMILSxwIMgiG9BZZHpT22DrpDajYcVGKYBhRwV+d9faiGJgJP1M4mJs4KwmSsjW2ujUsH20MjR
5OzHqMSTKWlaB4th0wqDhutMSuTa+a0PAhe9KLK1X8f18UOsGt5qOKy8EBC6X5YAkUCSps7OH29P
y9plHfCCKl0Z1wpWBFV/p1rRXNrOgREMJ42UQMYc//t4SQMCJ4WyyLYoxCFx5y0KN1It9sPlOBBU
Aqd3LumBUAio0jwNN2YXH+ynzyuqjfX4i/AwDKd3+qeBOVgaiFDwlfx4hISi+stBjBj2KEevxyDV
RINsM/LXWNR3O2uDsTunb5OjuIMyDCs9yGJz7itmwkRLf0M68Na/NECuYOpRGQOchRR7/SMSPmE/
qo4+phbHO7c7bBzGDMKAxzv0syocBkW5wraa9bNeJm82En1E+hdnftRrEq7n5CEn0p4dybxeuEYt
sbe0ZS+nQ/GkgorgaFN5vw4ktNntMSByMk6xxSjxsoniorBrmXuVvtd53meyyJlB9/HovrbTDH7W
/v05NTMu9NFqvxj0qNunQFSqVwSX1TNoNtgwWcghSi2DUW4UCkeEHiHBElylL2N9k/2RjhKPfz4i
XpeAOKRy36dN2DoYR4I+Aeifg6iemJmKEM16Nl60DT69cdZwUwHxpoUftNWefEm5YjKlEfpv5tRy
dMWJ56fh+i6Al9yoowpYDSCcmE6myp4WIod/O86SewtJpufm5ql9IIjFlkLhryw7dLIKJ3mDkXXt
t0Ga/Mjfm2RSVYb9WglwK3g/ZyHuR0iZoiaO5nzvOOtx92KbKe4U6lAshB/oRYAYroxarzqxtaAy
m8onkFZcyLP/0RUEHX3hUh8LgjElTPz2uP76s4LfPXf8BCWK5mn1gWulvR5yCk5wLtDGDiydWuw8
ycSO2Re5bd7YSSeWHsOo7YYVy5n4h1/D5TlVDi+pgMMErHz24rXDZGbrzuqxIBTn8tAidtm5NMsn
7pnh/IGCdy8SE0ruiId8j831nfLgh+QUkrkVPfWy5OyEWbNAUlkSP0ckU5e74FU93XmLBVQXM7bU
moCK52hnlt9KYnz4MUtWIwdr9Pk3AMeZpL8wSwqyIOSkZTg3HvbwL3haBLmvKNpo4Fi16NWZaY1W
8wlikPhf4KQjmXBzYEU0pErGul/0smeFWXzqeTMy3iHmvPZOmiiP7xBo9NnnxJszZp61ljfinHyh
rskigpGcdHS0Q/m2CRic0nzHxbOe0B13XXHPsErVMxbTCFWT88ccvSjKxjJQ8GWt9KlBqiSDKLRg
JCdQ4Kb1U7wfsH5IVGEoKOTwKG/3oYpUeUvk23OSuV67k9zFe11RRepxmTLhS34oQJfVl7OaATXU
YKzxu2LBHwrKgzgZwkt8M5BnoD4eH5kFkZ4QORcdD99zCEY3nWM/o1OYR+cJUP3oSE5azbexN9d1
jb0txItpdKaO3PJJGJR1ZOTR1woyBHJ1HFV/xgvHp20BsVWeflmbE765hoQ/KquzhkuuNJeHbeoE
i6lgshVZRcmUBAtU8j5ssUwhE3ymCEd32Lu4jdMR7yrdmu8TSAr69VTWZefTtrDb7v+k5orkoVsY
khgrHcZI3OLvhWJM8MTmsUEbdHnvh7u1JPw3iTULkLAXxrrXKX9gW7Utn8XiMx8kBh6N0buad/FI
DHvkDHTM62gdEICBZOzD2TryMdPpCFxv5g6bzQxvck1xWPgFcDcilwkHHtIfNG6PmCx9yeNRnXnY
SSUclF2K7YST6bUZruMkOetc1id5wg+w/+IwRTNQiqiHiOH7XBPCldNVaOQGgHIGqI3/UXYNVoqB
Ib2SGCBlBFvPUWnWmldjemIuFOCiycN18HIy0atLOcr5ysqwkB2mPdOvotRAIKj08ztHp9F9RLyO
oM/M0POkspOqs0Xdsv/Oqw6QMjikStPQNyxbBZY2anJGmekGfeMC73od0J3Sq+DQRPOmbklq5Hq6
tHhxFq84h9GRkGwFiyIvsSPK6Ufg36l11XxCzOxlTeEG+1aDufpC1Kv0URx4Itm6kEObKUzu8PeI
6k+HjurQMugQ1gCrM7JEGr22DquZIcSBkddh7MO4RbUFjezzWeu6nM4nSthZiRBJb4nnSy14L62/
p43BlQxOgW5ACt+5kKNsiibrU9EaMgclGF1czyKuKGZE0/KteP903WSud5dXzOF0YTmKMAUuCked
9rejC/DpvhymEXqF3XXXz8VxYqQZf78rDZ0+JdgWiXfcxXKuqKMx/t/OqC1j1lgN2kUv3iu8HRRb
IsaHnYNwP5sDz/0DzBB0bmxd1E2Eb4YPcAIxitI3SR1ijolQ6yrPh9FpKula3QQYgX2VBhq0dh1o
JSrbgs1dJn9NVRSo4zXYHDBVfdXnEWliralShY9Q4S6pj9y4JdqkRjuAydYHkSdfVOTFf9c+lKqI
zaaxJ1q/i1LzDPl2Tz75OwjaPFFtAHC2sB1VLmMMNMrqf+zlatrt3dV1gOVciiN0IvVrFyTB1E1f
+d4/APQnJAjWN/JWlqfqlrm8DtPXu0PVBnqCfyPMEkCpJazDd88oa3p/uL+lyJylY1JXLVLNrzhc
0YfIdm3Cx/YdhUApp76ZUX91uFuKyQMuA3btZsyjBvNgE0fXObx1LfEjc3o65miVreja+VVT3Txz
5O4tjtOnXC+fF9RQQqCFSc7NXWNbEyLhfl4OrQl+wbm7GZQ13e4pdDSaMhgR/twxUBWgck+r8JdC
omhoKo+D17Ejo4NfYX4SoS/ivA9ZJrmLyZF5/p4qjasiJnSjAARMgVTsQuM49XlIJT4m6EDH3yC2
JematIIqlezwDlrnkL66SqK/UImfsphs7EuRQ9FNbTSbFrxiTSazp/F0zhQLqBO+d55/aeJ4FXfo
MedtSrlabLassnlqhag0A3bCowWJZf1laNRz3GEtmOGMaEsBaXlKJhvvpbY0c5oLWGCV0Uw3ZCtb
ST3k5dqTwQLh0FOxsZLFV6ld9nOFqxpfRGJjN1hG8/UhuDjltwV3dw31EQ5MZ8h4N4eLAtk054nL
TI1MPgyG08FKhYHsvACdZx64GjjXQR4HDfG6D7Zdh7EA2NTrnl5dyORN9JkENId4A4OkvEfilcOT
hhhKwEoGPmSz7mE45FPA6IUwEUY90yB/TGGcQRvDE5fmzB4pA5wkk32PGHILyXc/OwK++2mVdnW3
Nepixa4Xs8uYHNMR8Lin/XslNV64sQCyRLFdOgTXRxuWv182lao8mttvItS72hhZTUXa02D/Yl+y
UzmyPn34LEiKXsD5FQ7bnIM5Hwu35iRL6ElQ5apuWktzW/JqjGxE7aSCnAly2W9tWsPI1ZAGDT//
oEL1YlbORgy49oJoTO6KKPdlIJkaDmFD7a6OUWWJzkMKc+zyoaE9k4ec6J1c1Zfu9gUVXqsipOhc
a9Noj1IXMIfNqhZDgGBgoE0EV55WB6RDF2pdqvJTBr2q7W+kyIGfRrVSSGpPbsNXhQGsy/cFTWwJ
CCGW9BIOrFYKsQ5UVuUOtciyJ3oWQ9kqiB8mayCuSh/JlSBexkzsKdP6Nm+z2wG235o0UzA64Jce
jbwdNKCIaS2T0Wnj0YhX4tF9r4EBpd6Zch8WrBhQkKNGwH/vZbOUqV5uM2KYLMA0daNmCjLbapl9
b2H3Zsy710SZhzWQhJ3PhpWpP4quYZeVLyA7PFoZDdgsShZG8aT3SABMKsr3V0QYbfVf47oX8gdR
gc4TCcgmjY1BsDoerL7YKaUI11Aq+jefmkBqaLfDcvPgc4YiBHry+KYk+GUQv9D3H7eNRla3fxD1
4/D84EpIuf++NTjLDxv9Rrq3xE+L4JYvGx7++bTWaKFcZlj+hbQ1pjZnGF6Q+cH5RjIZV7HIpNY0
qJnTFup07ChPl5+6tnpbxQFCIyioOBq/3ddDWZEb6gwtoGSEEFiZpsqF+1yDs4nDqdhzjh1MhE4W
QzpYHRMmNy4t8r4sumoNOmOLis1ijFpPxUeLVmLrdokaxMqHTVP2tf7CfcngWbvOj2nO0pVGhJts
RE3I86jFL01ZPTYJi7GWV1cM2R9iY4sUEL86ZvsPd8zO6VhkJUHje1TLUoEoDzRdJlWnUDYOIcF9
ndbdB4N6VPJnfq6mOp8Qpsl3E8ZRax/Bat+T8RgjNDYBouexZupTeL5QoeJ4Km/VdePAzTlkDoWx
T9u23IGgcY+bOspmJsPxRgYjuxxlO3OEY1bas2LOLt+Cd5NcJPUUgjyLkKBZizNJvPQwLK2Xzp7I
7jdrqQjB1tqxRkmRKbEAGjdoE1iPDpB1OoYiIoo75p+o2FQ0mhwcr87LENNY/kIri7zvrZAC7eaf
jzqu+FRk7IFdh3J7tpfE7nyY0WxJo+0pvWoGtcOvArBRIgjstDrF5d6uFX1vElQodyOktBKAW/lH
XL7Awy1AOI1gSs+8gdb8rvATUoRDkqm+5VDleREAS9b9nlhMIZWJp3qVYn8/LNU67fLS1MhakM50
OU4wpPkviYp4dqKfaYpj8BzJjv+3QzHQr9oPbAHVd9wfdPPUxAyLLhLFzmbhJJPi7h+BquJehUrd
x/jGNdTui+RvP/W0GfWwt+dfjvjThjvOW1J69I0xaqNHxcQ8GnIXAWWuN+HKuGzHVmncHgHDJmg4
jPnuzktyHxjEsA2hhiaT0VzQafS8+l4YVgLwzUW6dcsE4OY+Gy9cwNbnsHSX+wrWrTPmm90kVkVK
mTSuLmSchZjFGEjx9PgbLC2ectwJWmHHAN/xg4ApjXA20Hvcd4WmUauYX0TyyZScUYGyxi5dNCBX
AyrHssSRpQpM63ChQJA47iuFc/luRdApZBewElinIWIrwy7MvF0wGwDLOhN0dTg3ESlqW2K+pImX
llKU8j5JrxU2kdupiRS1oOnaOZjkZ0cEe1dgC7Va9O9Ewb6ZMcBDIpBrMLf6Gj1iA1yjUh8MZa18
CQAR0QXZykQvjd0oWbRwgtsATJbSp9Tv9M2JIZRNFmeFmuQrDgFupoYT5C3ZiQtKHnq2jV9vmMzp
MLQIN0Y8+I2ZN5jq8yKXOKuhxG00p+fBGWBOIQuhOGUA7CvGoCzf1822n1vY4CcA724cwNBWygHo
XxKybxChzR/HGaPmmWDiSZ3SHyFhapPhZaNHGHMOMeHhmw17KdAQF6yJq5co4AfVllor8xKhTpvk
k3TloLkX8kzrG5YmYXoZlq1rNGbJqPDpXaFhy9oyYLAz+S8h2FvdL8KIiLQsxawdMQp6YI+We+kk
QO7HtL+Q26zcAIleKRQPJATqayul++DtzPA98KB1v2qi+EEL2cr7d4LNUdUSkYuf2WZsExJoKOP+
BzVYP/XbdsyQNPKW0la15v4Rxez0vufDw2+oWZaBtL71kI6TRWg1+pNtREI15Q6KLV+wtRX5MDHP
TKj4jLDLxYfEYzwH5T9grn05pCsLptPgwyhYo29t8JyXL6u32ZxSDRqmxF2ZejQ9R8cS9I1wBCDh
bqMa94OQTw8s/tF5VD8uhEvSQtS1P/BnqNEO0262S97FP4H7e1mkXBDqWBsCUacCgYHDrsdFfHjJ
3HPhZMX8hFKB1sBWLlbDUr3mk0L0IZh1H1qDq/Sd1dNbfpx++YP8Zhqs+O34t3v9k0fisCm6tzbr
cluZYY50Q7YM4vuA4r2VnOfaIx5TqEQ8edSEGX+QFOl19pUqWk3vuLjL5yvhpThYJNHluuNSci1j
zhgPjj1K8Gh0/Wzkx0aAEZCTmQMYzKtFRaRF+FOIQCDVJ5Gb/u8X/GxT8+kyE6kzugacNezAjj2u
hoU6AIaNDKud9Q8DwzOrsE1SIEdi8OjM/L5LrH1IK91q+CCdClwUMH5WyR3gqie/KPflbpyJNyNn
32P1pw+iBGcGGDdPT6Hh/qtnc8y2lWu4DfHgCMluoAXCOscVMLrh3Ptk3FkeUO6tYqCz/yQit5Ba
CdpG/k8THjvu/x3xaJt37mKA2ZCfREpdWSJGasKJViEQ5qFAxnb0hbmO15zxlk/1ZEEDsKLwVQsx
UeP/khgEmqirp7HpCDPGFAVsmOXtvHne5Rck+U654XucgRhzm26mv9kbMGYUiz9EN+8uDd+n4tqS
zsx1XnAh6HGcLz6lPHcvMOCTttXNv6xgWUYBWAX1XzbVZccwxqTCxo6t7hoim5vZYi+BGCd0wXK0
2I15Giwe+Hzd9biob1CCX0usm1DW4I/DpqmnLg5u7TrVbTIa+2b/q6q+0n5G53qD0DKDKhU2B+NX
8BRMp26dPfU5LHyvFXhKe44a8Jl/BbVtD/Ji7W2XZtBXFJ+EiAdeR/G/3lQzF3q5fXsrRFJWvBiL
4XffNf/NsLJCU7liWS3h7CwC7cjAKdTvAxnIijx7J0KRRv6EGWQmDSvOaCsOrb71ibi2NTugD7wi
FYRbEdJvEOQ9MjE/+vyz30pqqlHybVhCEyrBLronpeh2QU4hRM4tBtvnadjMBlQV/Gg9EiLeLzL1
Fdy8smSDgIPxhfpoZefRJxa25y6DqSH1T2JnirLFkbey/m4d24CGEYx+HeQ3LADYTfj7gliMjEok
V8w8Gi3i6Aj/VZnrAuT+crGMwq5Ag39dlGYVZ7Wov720zgh5f7CO1cqwujtD2t70i158V829gV7w
OFarUwQoZIlBrVhCCw5jIDoeyHQc0Vpr43JGjDPgs8qep7OcvBhoTJ0d83NFuzTsXKpJ2GY9Arm4
Ih9ST544lzPDbM3fECVOy+AzLZiykh22LFEw+X6RG3js9XvuLkogqnS7MQlY9JZilMdMDqh6s+jp
QM8+9nXsxCArF0M5C8Tk6RWftAXqUfmue4nTkngc/881y8tdas0L598bqlNhZLqICYAUEjd4ClrL
bwMwIkBpOKV/RBXR+0dYvehvYM9yEE005f8l07sH4+pGJyoJPmpwHXa4mVIwmLA++ECvnXaI2wPF
780z7fpzhLiT1QjVgzxMkvur+qP4e8Dije5wZNQjnVX+rcU17MKnz8VaUQYZefY9FjEb7LAggtFP
WQD6KfCtnDAFWg+3aVvNqQ5Lcu6TR+PJTS+iA0Bgx62DtRUdZqdtfK1WV0W0008tL4BfqVoHeRQB
N/0WbOnTbmOALnQw62oFfUfFFneVER7xx/CKapChrVFD19F8z/YmquceUTvQWhjWFwEaBli67poP
z38zVcUT47rS6Z+fLictRN8iunC7vVzVkC0JsnGjfshYDR4P4xbPoQUOO1/hZsYwQqIO7RTlSDcp
3fNfqi6RKq6lMwo8SO8y7/C2pbCrjyTiN+U61NKX8sK4pT+a2ivebOdDua/6mhK37aN1QrVqGf/t
ctt1NZQsyRhQx8oJDC09BhOTgFbQ0eNJV4/sxKqAOhSWSbgd8E7+b5HphZOdK2WdnFevGtDI5P6x
ukQsqIjClq0VxIrr/Cyyhem+xKKKr3iW7Cd2D9FfinsywDqE41J+JOgNLcB9SlixK1tpiAbmyVbM
yKC8IvMAWQb4IsaaUYCUPPoloA3dqi+D6EsDTWTGXH6SbLDnBt6NSRVBr5olw7Z5WFWqQdOWpznu
P9eJ4u2wlkuRZxG2MiGQhrddPVElGc6Zo/ZvFZfBIfVovTJtph0EwtkiGoH7DJhmFnmebBD4Nij0
RwcGhcrEqufzh09ANeHul5K8QIG1vyhxFVQT6qr9xIWjG/DgAzXqcecExYzrNdKl6iQEC4vkdiMx
Tn8znU23YxZ4+tmVJvbkkYn15nFOHc0bBerkgeBUVnGbVVPJ68p9vsDAK3L92C39xlD0J56dPHHD
p34EinSP0VCKXefrxDkg6t5T/vKnobfTuURuEl+31qgy/iwLN96S8zfd4+KgJrBn7XdvWcfaws0m
yS2+LX95tC8wp0mgZg6R1S7/F7trNHio1MyuiAcaDNk9p7YbHaNnk00A8IyK2i+axe1oBYkiIJv3
1x/bg+6UZdFz2U+TdZdeKecqXW0y9IuzDE+yB9gH9Jvwndg/YSiz6LUiIrwfCOr1KpKLEdLdVmiP
bcDD10DKZetY5har+dXo/DbycOLPabPJutxsxs0O/0ol0o1L4wELcGnzc4k2ZderbkUE7KL9uS90
x5eKd+IgxW4zJzQ7SqWhDvQ0/LA0kTAEOBxV5PGhmjog4T0IoLJkXG0mnfgL/lnHUqM0L6feuReV
pKty85be+M7jnZ2QSwrOxHt7Cb/wxMdLq66UBg+6D9fj9v2TyAeZ6n0uEsghCwuBmJxyAS6ganoH
fx4zjGm2td3QraKjpnmaZYF+Td4nKK2hiDbvORyUdeo7KqeipF5AhU8IvAg+EEEV/JeTzsVAbnbp
/irLbN6pQfHpxHpzUS68TIvQInttY+jxDXWmpi3RmXVaNxMGvWF+Nz3n9AnhA5YH3j3i7C15EJoH
CO5mmBKQQusX108ggetnOg26zhjvhVnw8PkZYPdLXj+JXMW0/TAxElEcOWzvge5K09UTF3obdOnQ
i/CGRKSEMoCYutoTnzckCxccRIWACKCuYo33TP0Pg3NmCcMxrx3tKMBJHaCjmnLEZzAfWBFv7gnC
8D9lrUc4G6OSkUhd+qf9rBr60/HbV8tVulVob+IyRlVV527KxgIgA1bIDihIakPNAVfImGkeJzwv
E4lFL+ZsZXpwZ8eMn5UzMmhp7DZhjXonB3TpWpWa+SRE9/ysN3MICNbCDHTVKKW4tufhh5PzZokx
CVDXe4jbfXxx+tHNCOBiIA+tAMF1H1QHfm3EUPslo+roO0z5RR4TxM1ZZqYs3okZy7yxzBq6oHys
iLHRkTMgwpMMPt6ZTnJKvywW5hC7nxY+Q3ngDHrdcN5EPm0c09XfOH66MxXBKE9H0pB3x9AwVc33
C7F1qaMUhnTpU1AYwb/aRUofIAdqOaByuuDKqQG4lnKC97nCf7hrDbPquICIS28jpPruyj2L2cvT
Ghd8fAktUNoaZisqX8U28mOmZHuDnChutWSnODxCrVDG+9SKNUW7xnf5msoS3jcpfEs6aIXPdxyE
xXGxiug3HP3WA+8IBc6LwFhwgSFbfz4+qwFHK5E+B2Fccs1C2yQSSbmv2Cz8qzQ6ZeqFNzMM/Gli
o1HmvN+AGEvAcczIzr++O8o2loftZKVTnWDQ/0ER+uf2/GnCtBs78mtIJSwpiZY+FafrL8Lm+OxY
97cJirpyC0t3JDcUZrdeXxjaYWFpLb2NEsjDMBX1KQis6ettPDvhJAsDx4EZQo0rcu0kZzVLnKcx
Q9F061WuKNtNHsfL6b8adGAo3FXa+AXseR2fBIxGt+38qY5rgzazT0KFFnh8kT6TMje/wVaQsabH
VbI/fXpVQd5AZ5mFV1c9FJVZ7d2cJe1Lqtotfe+Exbt6j0WxmstDJ17qYqrDyYjYz6t8IUtUWCDi
MRckT7Qo6FA7rFzfkxoZBGeW/Vkpsp35YwiNMwBcBY0Jzfrir0hn6yqcWHMLxKWrLnV+u69PLhz1
N4fC40GYsBiCgKwtoKPnXkTDUYroXgIiXHFXi+Cg4ue/Os9xmucH03U1FnxoG0RgtZXd4JJ5AOLp
GYhx84DjY+RSeNIdCuIQjVnb5h7McpzL2CROBSjwjkvC1l88J0pXgshex2VlJQxru6WH8BUnEKj6
ugNUbX6+G0SxDpZzRUrZZN1XzcBxKfjcFLPzBS01gmQo58NVjlqYobGIkwVPGEUncUumRi56au2t
w65dzLfqjemCPdEeo3dTmO1M2FBwnBpzHAZ/Tj0IUtzilr5b0FgYEiCBhfkDrNwpfszKmgcUTZZB
7MAAp98CaJzpYi6ZS8TMbX2mjgvYWfwxI3BZB5+tCrDP8t0OCZLdaMWzjWi++tZZLVh+XzBuD1Fp
m2As4XZpktenCeURHdMuNWa7jFu1EuyLN9bTwxVvyg9kjyZ9+K/jB2UIjxMjAzqyacCOELa26TdL
gr8XGbAO//DbQD41zyg8EEuYSpcDdwhGCVNnT8tLaxBBDW8GV5gJ2O6B1QIkn2dD3uv9XQjNbBph
ZzsEqZtcJgxfDEUKhlK6AvPM/dRgcc7/G0QYNALSTJKDiA/Fdkg+YsuRhHLDvwA7M0gWEoHfcM4U
KRh+c/NTtH6PJqRwbuRNZeXsvyBNQP4q0Ri0Ys+LhGNbT57pBiPRZXBlCjuy62XGX7KsYVaRzco7
pzmQ7CptBp9OfvHQXGn9N10578zSQy970+2ZRLELplwpfyz9b//V/NTd1588N8g0OlE7xfZEsrg8
icsN5MhoCnafTjmmJJ0fdVCYt4XSVD4R0EzWHLihutFbNVqKgybkRXGW1i4YN6l1M+L/cjOCaaGK
cHY34qJBWH/nL40OdQyHpNl8JPd5JZgUIdBI4ZVwC5A37wvv/BnKwV2Wn2wZLGzrFZx66yYemx33
MPb/ndH+2rWg2FMnWdNHrUMvicsCHuiWRc2PuNnFnQEMutsYLcedjQz6BzMhsRCiEw/iB1+vCYyt
RwvbHK0lE1TjCQlGc5yMjYfoSwq2+pl98hsLPODjI/R14w6liEJMW4IfS+NOBC/iOA+69kG0uD2C
iua/TsspZpIZxIQeW6+utWVCPoqoV/Vn+DA7km8m8MYaiSXFaE43F4nxxvYM2MXCu2l8BkUq94ex
FX8stALaaArHR7xn/jwyVBdUqpjib79iBNwctP+L7bjENQ7X/d5HhjxDJt4zydFA13r38lD9ca0W
2Ufvpw+Ycflh7npdTjjFAN69Uk6fyg3n73HKs3XVA43UPjcICxiJ4cVyhmM7KyZnY+X9yNdkw8VH
eU9SBYoMGRpNNBRoVLZor9y8yqCZBiyKARp6MhG2bIIpydHkOmBWEVrijyWs3SGjcZd/bhIXQ03v
iFHXkZzImx1xKuK7npOMZueEvb+v138MAqUgPI1rrEZ4AvFVLs2wyMSO43OjfyLgg+wx7uxrSjgc
xbw2r5yyiBLuHxkERd1F/cSdbcj9kMbpWmd7lXoIB9RBD2KMAwq+eSp3h6W6JvdFdgSE3iak5y7D
bokNjmfIVwm3Wf3ge8RM/zIf61D5XuAZXJfMjR45FkMgh3FWLF+r5Uc8SSy2FHVoVc/2FtTRUhra
tXiwU2y/etLUEY9cldaiNDIsMzZwSu8hY3Yr9IlJ/diGPt99DFR59u4cTJmgmheKTsN4W+z7StOo
4i4ZxHXFMpK103mUaD8JTpn5l5PXJonVjycpZVK9uQvyxKv4DTuuIIzrJcUoVWa8UCo3i9P77zgP
RHJw9YMnV3lIS/r5HKKmCcHX4oBU1MnFlFflKUfAzdkWxe4RiJjxyDZ94597IKug0yn1YJO1Vvt+
MYlyf8FpPPeSV+W2QmOQHhNSw/wW9Aiq0oWPbzxF7VJ/LxGRm7bNH9jOQxMB3faCZpl8skiFPQzN
+5Y0TTi/xvYjRZ74jkGFSwUiXaMXKXpARMa32FQyNuuENRF39Fa0By/VrE/kSqwpm6T1AYnLJPhx
yaAI4I60eWsLd7cOWhLdfxJr9BnPxWuARxkcgZ4RxNIuL2+HlEob/EyyUhlyx83mVG0W4GMQpOSA
lIFYCFzlf73M/KzxrWaTJabnEz2tmHQpuN5MNcjzvj3KrEDBF6OjIOCq89Bx5mrl3wqw4aH849wW
64c+CLIV5K0WZZJ8NB2fJKVwaEOlvYqNeP73UDu2OT4SgDJvjVq9o7XV8uxs98/dmVtyrdjITerw
1VvChtGVY5/Mld6LXDiEDgnDIgsthFRQm6oldGgT6EuO5VuaaXqbKpz1txHufnZ6zvcHmiX/m5c/
OwojMulth0eeLL/KynFSmtiXM4BFo3L2EHgQfV5GQY7j2RuJdl6MbLLYdrY0xOaaAcJ/Al4x4tK/
1DUdHXvpxgnAZGnfvcBv+x+dAoTv8CrI0FTfb+qDj0Ub288cf6No4kS5GG3qyb5KpBsEH1NSLlHI
xfDhRfjqKjFPUWhCX4EEtAI6yHpVqUbNjS5fMG07+s29CVjGhB3DyRSVkk+uq4hYAWhI859ikI69
0t1NASpywK/nWPgV+PIUCy8iPs3TY3hN4cwBrXYEVAiVUDCkl0xY8dL32N1EeA+hvAxD/lqaI3xq
XB4do/YJRZszzltulQWLNjYg026tN+vrS3FvaFSZUpO+ZSQ40wEcG92sJCxDflIWwyiCC0GicZco
A4yPOxtuA6zvo4+GMINMs+l5VSo1NsX9h+pMZ0P/AyTwUopzbvhzcjqIVmcR1P13W4C3Avhbx2pl
M0rCGpFlB6YYtVKyiCdFoDGOUyxe6VRV5S0Hx7Nb5sD1aSYAUBrPtiA57J99ZcqoAhlJTRNows7/
N7eZnW9f+FoV/+VHePN7tNeUL3YYSqvIS3nfG9jXx1/hP6fERXoWOoAl96yMnck4hei8Cdwobn7p
7TkXEQJYQpq0I2Hedll4nP5GkV6CiiFqtkC7/Baa9vnj+ZWL84mvXh7KElF8hweJIIG+pMhD4G++
/jjJY1NFhs3D9sj9okpGbur8PURSLba8xqcv4tsiauLgMT1N/n2m7D2GuvJF617bSC1pwjrJZJXm
HQEoMdyHjDEIMQ7PVF/vXYq2wp5D24lASAcrAxQJsESStlDRi3/ipMztoOMdy80LI+Tj6alqf+sh
8hVfzJwzR8sZNxSvzw7Lo//QmcyP0RyOsDpNywLQqhUNUA3vCBWyJh9tcAYIop9kR8cphuXTX/Q9
l5jBSoRDR4GAI4OkgVZmACRoJeu+6gOtCnLkgJuGp5fCIKdZzyuM5yZ4rNvhXw2ySc6b6eYlUjYL
lXaN1TrA3HiyLpGyJzQyNIbsHTsUTYQ0LjCz9acp/BLflJ7NZegy7OVh07OrCkUI48awcNDomjXN
rMUz2EUZE3P92duXIEkrctMWotvMarVu534dCx+hqjYmFDWDtrbNWSUq/ubkg6xcmgtIcsPu/JCB
QV3soGsi86rDTVk3AHVRFD9Do6x5SOpH6E3TdpVh7vDrOKccpOmDFv7reNF61DZ824JALRR3dMWV
q4L4HMnq4mOHWFMLCzHENaL2HB4w+sfUzPYgRM73/67B9XRJF1Y06EWHAJVWxWDs2U02rM4qM8mi
wKsDF3fVfzas6ruP8b5eL/SaOGEvKmR+WuvuKVcF1o706lC9Mu3TxFoauCQ8cCbx5BthKZONjS+n
hIJbwQJoXDb+cd0zIEzpXINBW6sF6Kmd/LwQG6r5ritVclj6CuTBC0gJH8WrOJZM54VFJsaRf5ub
L9mrB8mSzSYx3gOgG5tL/h2lL8gSpwkC6gqBhcAObNZTgk1BvtKUovr1iWF/b6Poyg7C9gBOlbJN
SY2oQt64Hi3B9ClSusmponWc14ZhKne/TbzpxOikaI52mlbXqAFTFrOHVi4EE2HCdbrxQDObs0Gb
N5CPzp3z6y8R/ZaCJ5L0My+QoxOIrGqI0EwgZrgNjQWXFm0Jpz0Ag1VDHvl5ZF6h3fgMdSaP7IIG
OYuYLY+ohtytk0pMVBBQf+YPAYKLH11jFrgM6ttu7or7cvM8rgQKQVpjQBpQiuI0J3UgX76EAstH
c5CtWkHuiTUiEQnCfWwBE5Gf4eU3QsXCAH4vWWAwUmSC2PVr5u7nXfB2GbCyxqyPHh9MlP6PUXFG
uUJzfWbxSELGjoDNdz6B5zf6sxQL2AHv2gkjHe47HQtvtVRBWYDeLrHgx+yRUqhrLKbIo2Oyk8hY
7Ffl/3ZX2slxggZhXAHSWtfARaiLjz4PN7oXV74EabC5WU3ebFtKcKFdRN7WAbanOooNf1jAmD9B
lRTT2jnz7G48nKGkOJRFvXO/fhwWSJjLKITUn2Y4JJnxVObJx2CnCfNAG4akKUXtTdg20XRrRebB
pFZsXiSguMqcCnBCoX8kms245qxWCpVZxGhdzHlHT2SA2pHp3fnrruakobbA1Xz3Xj9thsnQWGIE
pGR9NOKYhkDZhyKKNsQoywaUujAJRIeF5vvk69mTcRcT37bqjWYxZdsSLW5e59ozdbDArVPLi8X5
a5gi/ywHighEeVriE/oqn01QukUJ/l3cGIZRqcIP9grAyYtU8bJYhNYcUQFrQCj6u6XkU1nrrGNS
tmtjftmDJ1J45xr3erMfYHGFrgp2UdYWRd7a+1+pEonEqxGd5tOvV5MvYJO+tEQRfTkjNEUq9/vo
pTWol/xhuSEGVfol43fM2Lo7iEPaqDvMuWAP61DRfxp+yn5Qs0pEyif0qpJRa/Mkm7kfT9xvseu2
ERyD+6TNdVoYY3RcCZcT8rZ/aA6ii8LWkrNgBshBBcbPNW22YzrRmHIezDCNvP9ydzUWuQZ/9fPG
wa9/lrdbdVc63TufedvsLEkjZO2F+CFH/bPzQMVA8uBNNQAqjOxmTD5gs2opf6Ow5HYjXxtlP3N1
jf88SlqabfajnWJpV1786+R4cClQpGkrzma57sgMzEtIQ9BLzzIpYjBrzCayNBt4CIPKMrdMUY7S
zdQ0kg7SOKl+M+hPoODSyy31D/BxIcx1Jd5Ke82lbvtUbsdy2ZxGmtEc9N+52Q7l87iWA3TQypFV
9IJ6W8ZJLdf1E6HkG/apaAL8lZOdqXzlfkhyuM6gDh8xVoh6e4jqLgPaPO7XNUmAOjX8os2fexpH
nhtxUCF3AUNnNxMh+5ssomH+TgTYWB7gRL7Q3X2+DLsWo6seGBmYOaWOhJQwpQZaxAyk3zImtOOn
QmuK0VynlTdPWAOIoG3xc3HRb/RAvTd6rRlSuMKsl5N2GNpJBqFz4V7p9ntdQMphEetJh+dDJnE2
k2e6rCa/bpfpaOOP9Jjr1p8+bkdsz4dRCsZgdaasHA2TdAm5ndrG+SReZE26E/iSSeqVe2hxroaX
VeTLSYVEyvk7aaPgxm5fP2fzm2pvRR9giIR0ieHNioAv17+ceUfTPitASNGrHOGolQ+cUSFi4f1e
N9esGrQg13D+ZpZL31audQRkw3dhnGEExOLwmYXxjKK+c9HlpWFYGwKXLKRTYSn24ZwgDdskiF/U
3a4HGLBbfJoZ/POJv0fI9+4sIuCwZwL6/qICUH86eldrAZFk0afrojuZNcWHap/8WzPzN6G4Jf1n
M9iTtHvv4Jqp4JHyyGC+dGfNXkN3EbBsf1La1DEe7a0eXqPyOEDDX5uAq8OA+uUCyjyuB8cplqts
tUUxGIc73GQu0sZeMHoCuZTktgWfGIZRUATmze4ERFOPWx/vlgQ2iqoGf6iyBIHhmm32G19+ZCoC
GbfZq9Z53UaNQ8eBuIv/bsRAvii+lvv8xk3bNbMRYUq/X9EfLynvPOGTRPpGkj0n99TIq4d/5oZ6
fcSwkfHX5yarvPhkqzESfRp3T7UlzOiYfpZa65aOxqg02jkxTlW6VbKr3G2jGa7dMQGjJB5glv5u
c5Qys8rofhX8cIyfg0RjzjgpZFzyGGaWgS6jwt01TXoAh9TC4C9N5GZJ0HhBx2HrezV212VBmiyW
MQTioAMy+4jM/8do/rQu8Gl38RMplNpzWen6vFjlypffZ7zAuzkEQIbFkAjQIEfc+Ol7HsVtVSFO
PQT0b3v9Mcj6sH9n4eJB3tJg4F0s4mXjPSOMUZ7bFEq4b7nryhJy4fX9lLns6y0mW08/qlmJM+WQ
eGYXpSOFOV3FRoEa56Ae0cKeZtXbvRZFzO6jaF7P5700KnaalftQ49aQjfGUMFIOtWUq9QhrlMXI
//5VsXPORnXt4EBIMEySm58bLjvJu1lqyG1zKAetCp1ZUkXTHyOcmO+5UJR6QFcxJBmhPVNEBv1x
7/gXwwO9Lua5nmXjTw5rOrnidR5XXdAK86LA6FokYGy46bEKjnE+GnhP0DgNS5TNj17ho2yuxXQ2
YgLKjLFmy1Rgd5y2LoCYYAW313S4k61U8GDm4hPi6Xqn7tZjxCn6XzZ3J6WgwlBXXzt4nYWREMW2
VmydO3aOsMnHb7s4ZeMYHlonenZNDeyvf+Lkgtf36s736PoBrIlryBdN7iVBLv4PRT4i32e4ybj/
OKR3aCTIeANxOVuFUz1uCdConTwzWE7CzEYsZy/xebWzBO81jqUEb3eQTU3ArscF1JUFoDzTcdqJ
WJF6NW++iDb+jlt0PEYc/7VJ+OFdWkGPjkfr3CHXvQ8xgux6nmXPRZh4/5D2+KuiQLKg77eo72y0
U3P4Gzd6cV3LF4T6AQEOoskEKlIKdwPzEJFm769TwsS6PnqY7RqEP5/yb5O2ZNoHKU2AD+3LboxH
xZk6eSrBO4CmV6tjX7KJQwadbZCi2dZdwsx/k9x6utQedsHbuBIJaaB8reZ3AkcH7XrpjdnK2GdK
9pSQ8KBHqUNz88S3BAJJSYsN8EB+nULyYerkWvrUmNWgGV/m2RAW3ez71KnbH2uQdJNam4iNmfpU
YTiuSh+59v+aP70Qx21AEmgy6rrgMPDoVoUdPEgyQ7VxQkfKaFhSlm3XYM9duXZEsEVEMlWC2QvA
gr22fzvE+2sQqRRhknijVi6GlllrAouEl4f2tknCyNYPkxBvSDKGi+QyU7NmTZB9hwGFHrQQJVx0
tJOA9UJLyMEna5POqxCpoXrs5SneZGpjWmv0s1AzjCZbxbUYhGqJG54mO92j565Xbbf8EbSFHZZX
7i/5lnTkcQi80o/TcZfiJzvO6edLhuVcfqWo/QZW+p8Erl6/Jn+5arufx8Nh8y0r8FVVipot0YR1
chwELmHDGVZPW3EYhnXKH85502YFP4FERfV2eNVVN4j69aBt4oCNqJsUtyd+1CBxNQdK0JSnF/pZ
Ky0jvPkNwYIiuZ42441aZGt8sMMpm9PcWXOXhJs7FNpfWgyQJOjaaMHrcxr+NRHxnA5Z/6ng+1s7
5bHOn80ZhvgAPk83VjKRQEnHfp8oOc1FyyF+DohVvZaSCLYxKQNGs8zSWPBWoMx2hdSpFa/ejujC
z/z1peJ1mqn5+APklGVmjnno7iRcnqvcBvCKtPss24EIqUXWOtSSCdB6vfNacjTdKPSX2MTnPxao
6vScHycxrKQDpFuzViog3zelDQtu4onAfJdPIWNs0hPzFWN1W9yTGxu0O9NSCcrFKfm44MEU146X
V+vnc2YnVVkXYEV4ss6zytdZLKvAHV3gB1V91+vN6ySUo7X4w6gXcCCHXwoTxl9Zy5eZhe1LneXa
IL4hqi5ODk8Cn91rokHGCqBXV/QuPbWHe0cV0oKbRJCF5Fdn/yPSAUYPBM6aUeQw9MQez7dauwTk
UQPrPw3MdSJ+gWzKV2qAn3IC5cHsO9z5/6zzOPBctA+DvjU2/quTB0He3wnkhk0zjrVP0oN6V7MA
fir67SoBNZndH//nv6hVZUXdOY2WjpdLyGHxSjoi1xGLOGUztePFyhxqJXJ3RGExdgfdwesFJjXu
pSpSeoDYba0ow40CySdYQHKoH/+7wlf5oOIVtndky2QShu6CB/kW35p+CXa/d6g2Wl7oW3MItj+X
NLdqZTpozHgIWFY0+sr42EshEDFCIWqcNwFvDRUgKrFToeKPLdbhuHo6MZoxV5R1qrBsdnRzbIXJ
1EcOlXhfJYWpZ8YWT/T6TrpFpCvkSWkmSGF10Qr0OLQeNEk16PYv6mA+5IwRF4pKQ8m/5o05eZCU
YRqBsrcvcv/S+mvx6/93QW5zUT2moPTQYKB4bA55DMC/+C4+87lTnd8HK+NpA1IAfJp2gpfM3Ugq
H6LHz7o/U3xQuW9bsiKAYteq87+5Twft+4T3QQXykRNN5XEEUo+G2e2BP7rp9BYBqaGSXL+gz14o
pF6V4+26iW2IBBz5fkbgSQ4VHuWfVEZ5Z9It11i3VGspbCFaWJcDqGirRwcyPDhibOmIntp/OcmL
bjhT6PxCsvpsfHRVOPeNfQZMttfI3aEI+o+bH6aHqLC8H+QDd4fcI9uuhTO/QPOOid7rmJbmzAzY
IROzAvnOKSUASNgx0LXZkRbQmi5h1FaEBSUoHH0Gom80nVbfcw2n+XdaZ4HiCspdYo8cF11wzBq2
Maz39EgGE6BHsGMMwK7J6fbSqGD9Ndy9Qzpbtk9vextIlX8fWeO173zcVBIQMtsNi4yH+DwvTfu3
EsSnUMkQFnfD0zs7eoqwx1xYT/27Pm+cZyxtLk2X3SO8n/7gsRHmn+VzeSHyIs0xUnIV+j95tuLt
pMfwhPzFX03xQ7XuIn5GAx3KndSizcc01SfSjgD/Md27BrkPjKWdIS1jhNsJTC6eGuNxo5wsX3K4
FWs+4JhYmZ9QpyAXtVFOEgkMN911oozUrj20qROz6hqVb+687fF3+dOiEw58POlWOfdInhOCMLRN
1skFNOpj9Ks2jOkGuc+Il3jA2xaMUdbWQY6s+DbWID0a91hMOzNnuspGM+a0lqG9hxC+ubEgIxgz
DFAnoxmbuByHYnEwg4TKmmZjWZeFqK+JV2IsxJhPGG2F8VhHZyQiPVKrFcW696qZ4QCKrZXGR0h6
Dz52EI3r4ExTUr9eoXrcGhlD3QeaX1sTE7IaF73Kx20CkI/nxcNk2aYIARQ/hYgbRVsnrShShU96
ya57GRemu1xCBPKV8nBUbVvb1jEKmhbSIJbvkrva/EEXhkZUj/1Ld0Rf1utCQ2ih6Q6LmMyGvpno
yM9t6T51tlPl3MTT2sGpdWVqCL4QXkOzO5ykeDYLVuP/szBJ5L3wN+QQBnvekp9scK6AawREh6am
1YGuTGm7/2MRqU/mFzq6j2H2Z8lc4wYT+LXaUcW2e1bErRnGaDmqw9rKm2XC0R7I4yuUW+s99WeE
nt9e+pyE/zve6VHK4dGRdoxHBixFXOs1t0qtjC69DygZA9WO3K2Ta9ZaxiuLlm4oDwh/q9/MWmn/
xuzkEX7LrDUwXs2fL/DTI4SIWU3+cXsTDDr2Clat6jpfs8g9XvPctBpy1iar0OI0SKoJvFdyzwen
vaCCQmb1QKGqZu95v2BMIZzV1FJXHXyH1Yu7ZsWPU/gMZLJlo8dwUywNffSegQlt+HZK3fYbKzQi
vJOwkSfjUF95zRCR4dJoNF8LHtxf847WT/Nwcdg2jDBY3tj9UmuIl+QE4hjBiAkhMJLkx96nOjXE
3plxnsI7EQo3Yd9vhQZzuXLDSorwnoqnU9nNPaqUKo3hWHQ+06Y2j3HB4P5pwsVB1ObN8TobCXuv
TwcyQ+secel7/SONVycz1A2CO5Nm/IIB/9/DCM9NMhj0TvPjULq5wKZO8IoCHgQvO4LuNWrnnTUM
Lm2krvZ+XSYShYNr9lI/BppcbXTulTWEjKcf0IXk2DPkYjJNzb1gdVulR6OwKem875hMMSXgusag
ol6I3C0ULdv+GA+fDOpUwxh05MXsEmlkq404MSKZY9USha5FflW3Ys2DTWz2can2FSxrQJ7hxW/Q
lP0X04nErukaW5OFd0m53PNNZceibvFpOysxrSlHjnJU/3DiZJvvTuHbprT7PWK17YuLi+FG1Til
5hgRpl9qZ2DQiWnfxJGQtasKvVm/p9Qh4F5GSEeE+RjIngB1IFRVjwNgQ/FR6HrCEXhTYPK83/MM
+1jykHVSZenV2kwr1cZvrNgN/HAgnZ3ZcUoE4s/tI6FA7vS6dwJk3Yn/hn8zv5XtUzWyTj1XBCtU
LFET53w5tiZyN8u04HpSB1HfscAG02ZG4na+yxDJKlqLO95yNQ8oZHDCrHMxt8GHyZ4fhqRd73/v
Fe6yN6Vj/BetYwyq8ZMiicV7HkSkQou4P8g3JiUmy7y/nKNfJiiBGAy2CborZPNioER+Zs4ACHdF
OZIAdgf1lnF706zUH5uXsMNBYw+XW184QBmPiMBQEBA4lpj2kzDYgocp0IFftw8SsBYF6uMps1IZ
doa8SWmZRBN5fNTPLfuRtYtFNIMRz671bkhBvv/dexglpfigSxoFXQVFYAPTsIpCIliw9SofERwA
Vw4JwtI5Vv6BXpJwrxdD7uD1p6F9HHNonUE83Wq9pTHcQQSFABqY+MbwC7bvUCJOIBwUvCu5SnFb
hMIFmxTK1lBGsZMjl8EGYAxPj/5KhQXFoIL8UbYJkmi5RUT5DJXspjYcIK0egUzlQbXSAoI/pQu4
R1JNecEHQROAruMD42BXHII7pu6I84UbmE30f6JrOzP5YlTpcnJU8smf8I5A5rPTH9CVr5JVW3rg
594a8SnQKNX+Es/XoKVYDCqXK3b7yMAiLAU2UAgVn7L1ubiO6OK+0LZmutHI2fzaaBb+70IHD7dJ
wqGW6QbF1CqyQGv5VAXanyFIcEYuZf2OmcNjbcCWXb3Q7eaLtwEUOm5Rn4XvRlBDkD0G1jDhoApI
JMWEDdq/XRYCstEWfRHGsyDBodfslNVkG+a5hwi4MovqMTnMvoS3/j3+cCGSioMsQ3rbmv76Bk8j
tgLl3UXMGAXPTmadScN0hXpjyQa83nEh9AEpJ3mK3QoCrODET6j2kDQO97PhhY7kFGwFzbBI/zJ8
xxEJNtwqgfm3pQtUQRnwU5oJD45FO4cVzf7DuKB76r3cYgKDU38PG2fFVuphmlV2KE7/lGQRHw+5
imXBBHQJg/LW6bAhiU4UDCnXK/193XO8CO2B1HWgWAD30zZqdKogWd9SarJNCr7eChs9RI1QHNO3
EnygR8DnnXX7K3DEJbaesJILpJ8FFB0gud7l6wmEVzWZi/Po/eeQZZTc0FxUFfQHTfR+HLwSEcL3
X1odgvwFMoN48KmVyeuZLkrxMtEsKtGniGOZRWa6ivsSYWCW66ApX8RhzULx0IJ44UROXplYA+lM
e/C3osp144oAvfWz11l4+EcUB+NdR54SUSWrPYV5vvvDj0Rd3Fk4xPEhpNwDVNooPWOlIefZv9vE
ROkb/V2sP5xXPxKIXieyKJJhjV5LsURWraEaJR6/BHXuLPOucudN+eaWCddIz8o5z8zZqIHPG1ut
xvABl9FBPatcn87b0TnZqBOxBDyG3WtrHvWkEKb39rHgqHkwhdi/90ctXk2Tgo2oQUI7OeBEenNS
MPLPo20XIRNQ9P1ylDpz71RE3+zT40vgKMs1vDDB9Xbgx3ZXO1OsoQHeI7kPsfzXabItXInFkKuF
jQuDo2301lfZbmlnqa85F/4dyi5DPQgPZYBNMQ5Pk4TKWTAjPWO/yE3cn65gBRMsj5Izx2tEFAVt
HWK+GEdoO5BMfVUFHvplsn/UxlA7109p/j5vaR6tpVxMx6mJ3Njrbnm0E+dbmqcxTbf+sjNhcN/l
J+JTAGG45MsX9d1FtObDKzyu/9E70qh00KvaIqXXMYVjpm+AwVdq0VbyEDzbvyx5mJAjoKRZGHcY
SPPlOVpWUNsLa78B9IMAYJU1g+NnM8pv+zoKdJ+B9uEC+MABNm0R55AJ/19SoojsvGk8+Ky9chEp
O/ncFT1bn14d6XxjRzvA43/YVlNl4tMK6ykY5FfFZP7usBVcgzQh7b3jPT7akWaaiN/exlH484b6
mZhkkzvXqrJzJWmquDn0aTDH4bqI92oh7Z6fi+pxy9YV4lQQomhe2PbUzDaBDAzzwMeaSUBGlpX9
L5E1RRZpVKcGdHtO6y4PV5001uXvaYdKiSh7ywsU2MT8Zs+Ld30FXa3l0yDW5pyRQPXs4lHIBUeF
6wjGd5T9TQw3alm4Wqf6cL9fsJZDTUFC6YN7NhPXaM3xPEpwHonGLfxsiglae3go9oDTL+h8cZm8
01wGw1udNIlfps4jNzZ/ReTCoDKUWCUPGuUcP9On0v5Kx/wrpfoiN/gdrbBGmEeAGJWr8z+WTUO+
OHAdG1QEMbDgm+DisNjZ2Uj6zk3wIBBWx+laOR0SvVMgzHn4wBB0aBEBZqPNmUW3RZgVvZoUz/Co
Qx5HOKiPTbdj0pj+3x+ML8nVr+NneIBbzhJhwiQwCfish6dHxUooRk+Ko4BNQxHzn6VBqx+5Lat9
9urV5uYG8381/+w3voc6ETiVYIRNzZcgNs7MyDaVhXSN2nMLLUeMVzxMybYF9MU+NB6mvTP2Twhb
jOGscvIHNmxkKDNTRdic4ELJgH/BDJ6j1sQD1Ue9/A7DR/BuklT8TrIq447Qsb4cIc8vqbxicavK
mI0ucI6AlLua0EjLQhbMz6bXbkw0g2NW7YCq6If5RefZz4JYVomAhkb316cFuXZKrWa4t6lg6mu9
OgYqwfGXNU5L6Fd7+P0OBt5BgvsKE1sd8b99tpvWraTZPRJuc0q5H6oITOQKjBe25tOKJxBozgGG
C0gnLO6qnL8UDnYbKkHpGps4o5ZEvlG8vq4ij7RS02a6ksBhpmI8UVpMn72gHjGK5D4MCL9ed47e
rhwpzqUOMBi9+emfmaSAqaX0V4cXlk6g6fGk0Z5Ryc1s1mnfug+mWNeI6KMgcvFmVpsIFEEri2RN
jeunMYnph5O7zR51Jkb4XCk2BdFknPkWSmIQHmG5A4zfFuptkYlKggnFDa24IcLFfTSss31uE/oh
vTULuG6nUmcM4bPFI3IWJiCa2zxZqLCjTOLplzkwto2fVzE0+BkvRtVtU1Rp1ozxPBbVp47IYAea
BmQo7QwAPpQ2CJOkAIWUn0j/XpB3hqQaCcd3ldctKE1fIg/PTcHTZCwCvIj3kTbRiaBnZ+4GBEZW
bEsFdSIocyskxEhD6NJOGmIQ+T2iC09x0hizc8NS3cDexBFaO3YvUcFcQkVKbNY9LDz2EQIUsF9J
TTly5IrE8WQbOWqbU8LzqJId3+v+BxfOVoCXrCFbqv4E8Im7pJEc2akT85TyWAwnGs9tbmAloW9I
O29e00tahszpkCn+Ov04liHugq65CmyC9k5g0B/bePI54YyGlNAZsQ4b++51vy63nyO6lDHqBgHl
onW/9wDx/O17nK6dsQxn62cP/eTceSz1B2eDSIoT79kfT2zMQe0lMPPR3JQKbG4BQTxQfYRbq8VZ
G5rQXtF2zih55mLZrtJcft9pGEpNax8BjHRhj0fckZqgzAmgVURNLpLCjO+IUANb9EfqR6nh0iDR
FXOsoqy5Wkq7kM44jI07OmjR4or9w2WFObNKf8AFkMDYXdVsdV0o2+4mN4QQqNYLg1RULDmWlMpD
PqARfZYGWSyPgx3n/FaarqY3fDFm6w7D870njBAaB3SHAZ/SDL2WLJCgYuaHq3i5/vbTMsEMLpPI
GSTzbuddXtaC3zjK8Dx1hRyLX0VrUf6QWl/G7sZ2a1Sp+pZf7bE2Zyu6v00lPG7OcFWUWVQ93zVB
xDBBzBx61M+GQb/CmDEZyDo76hFcBeXLraTHiafaBOhiWCuyNtqThbRNYKGqLRPeFA0BihBpe7rV
+ZA3UW3uOvIFyrRoLpMHK/ARQculhYFzqVqnKlea8oPwespfJZsctVvxSWsMj3RgDDiUvc1iEuTm
ck/ayOF/v5n0GHgXs0ADunrCm9TRzrhTrzSG6veIIiKTmm/A7nM+XoDwvT3k+rAWCAnLAMbyZNuX
YOPFd0ykLZEXc142WlLahtttSA+UgtBYx4aFgqhrNEtkUubrMsEfYpgX//9dvEAPz4ZmDKINGf8u
1qnY1cdf4YcabOiCBz9U0KIUXk/RPcrbgaBX5nc9bF72zUBRxU8VbHJc+jaqMsNdSpkCG9pNfBh8
KbKBx6nHXh+EDlgBsZZjZ1tKGh1+BfyGO9j590KqWkojF7u5Qha9H89HOyQrUmQe9SQ6wt4f4vAq
n4vt6YpliDUGiAQljv3zAps0qOCbLB5QDkiOu/GppGGx1/+pSG4twWG8iSm5uygY0KEyNBkb+YDy
+lUJFNC/dfhafz0ABAgo6BhG/eDvpcy5VZzffQihfmnmztaoQAmkCHPMAGieyHbMiT+iK341KED8
4ffY0muYlu4yHspp78+/xTmzlNiI+LtvctAEPzKnySRkJADJyRfcojVqHQ/1bp9UjKhvc43YwU2p
+2/QF0dzIXzduasouUCBYBxgnzBjCzUjv8QqSROH1aJxBlWKtGL/+sdz+8OEdOnPP+zqtkuivoRy
PkxgTl9EyavExnBdn/u/BVWSukqQoOBICj3kekvFTQ0DPChuuvsO0SSAUADHKqA33AbEUmgZSQLF
zSD6QFn2wCCn5yJ8iZt6vdqkE6g2MfjXxnnV7ENmP9Eex1m+AVNMeH/5NCuKk9llXtPqz3M/AG2i
y7pezATZSlEMDaot8pZHtxF7LnpFYUOPYE5drbD6WfNhUAGWRNFdCnkEyV5It6YI8+EYQ2gDZwfN
xBSRHkIMknMrsTT0gGic5rnNw/n5iREoOpwRNpcMoE2Drq4nsp1mQNzYaY7JlI0uavz1taWpIhKM
HblIddWrA2UQgwZxkHOIr+telV2H4Hw3cZYIZYZ/Q1MGonEeAcDkd0QIDmsDcDu6YgSNgQSrERTy
R/8sDHwnK+VPmPhwMRx5Hqj2Wwe+TOkF/DFhDalrnD8aoJU7f6uojfmA8NJo1P1tV8uR2UDeEGhY
Er0w4O44wcU9uBBEIMh5dTygVexrFw1OQeIObTnC/xIxhP5Ee0veC2yQ6Qyid40/z96xH+IgISxy
DFgmNOOTwnOvBJ/bJCTN6Q9lzcm0xX2lnpbHsyx/JtNohtlMaVhqSd4dU4sXZSQwZsVcpBysd3uv
TrWo8qod5+xs1hQZDAGjf7EU3U1B6vcsv7sbg1VF1uS4xQOLb+xxo+73gR3R5uQiMl99ijEeBnm/
Tj3Z37TQLNX3KTa7zpqj3gYpA6p2mTYLuOdzAEwSW7jvogDwUXN+qsvC1lV/y5cv+zIx82EdOs/1
9xXeRP7xwcwP8dxkqURGFQTVQ+KoRnLZSVCUKvosbpjCQ6qshuCBdsCapCOH2nz3lQY1EsxMwT5V
zI/KUsGtueDlxg2bD1TWoNOjooSSyxaPZS5G9QhLmlc8sV7m3zuyxtiCqEm28Pzl6xot1bY7XeSs
hj+qIKWCto5QV4Anw/nLPzUwxNksXrPWE5P0aNk+3ltpi9Jq3gtgK59p284JtLufU7uypFfKZoiu
oh91ioYtviDWguemGTM81ySvO8wZuG+c+1Ofp4pg1EtLG+3w/aslMXXX923XRgfJtqVC6H2PsMzd
0QXxaSJrEDdJCIieFZNciu1NPbht9VO3NqI83JH0y/E9K0+9zXFqLg7pP80xLNjP5KdeRadCOLyu
jnY/hNyJE6rG7l77JMwfV5loy4qrkjxBZjgGo6dExzr5CiczcmRZ+5QXT1WZjY6xT2htdP+oIiS1
rpMujH4kx3Wc5R6KHqYbE+8ESb2IiDSGFFVXIMKviuv0oTtbUk9Lv98imAaORuzXdJWcEgQY3Ayt
4IKBeSAv9FNKe6u3me+QA3DRP2GQWv30mLfr73vvJIEt9dtKYhPtyRW0IEE8DrEGNXShl6HvISVb
6NfQpUJJ4T9UX6DYHruKVMe5USQJ7nMAnuhYka1uQTUzf5iC9p1F/ea+1YEa2JJbQ1KIDT1fbOIf
bQfKT3NtDkCD3g5Xos+3JzrVMR0p9aj/LSrjkwwgn1eCVCNnFd1kvkB4vifUbjw0LqFC3STr3Yjw
GChpUEnDnRlflFfxH5Gn7voLJhBuD3r6QLizdCk7RI31ZY/Q/1JewtTZjlRFHoU0w2BGdyqDmpBE
o2pEtxssv0AI/iuL+1d72+H0R8YQQY1dD9wIoeFfwi4+qn99wwa6peMlgEDpbV6zVdyDlnAVhyVy
gJ7dov+WPz1zafAUHgKyl7hPonOww1x4jRXDvzXn7RKfzPxefYXfLhm9dI7dLEpF3ViNc/feVdhW
w5PaFzog9Yvc2rEhHL7hjYQoLKBgydw6krnMIAkBiDJiwAjlYNuiY33qWIbSS2ZoSdUo2he69m4q
8KP9Jc4gET1xXFerAFDDaJaVwOkOzo0vx8N8TUo5fUMHQbiaSdSZXNVBEA4au2bO/QmctHvvpEhB
mIU/MWQy2qXkm6gjdgw28mn1N8+6NbuXOLaeTY7V4McFjYr32MOPFwvuKI2lecYUmQlaHEEGZmsT
GMQfJcFFCKgCgwhnihYqKQRwUMV4Qfbt0F3aWAHJTJ892nM31VVmAAiPUxD3JynaLGuMswUWh6gr
moz/IfL3awhY1jCvYObyCzWQxvzxTccDuSulMraEb/X/Etdgd10v6N77yMpU9ipVpQ669eYcMGf2
oal+IHJbWgyLjVrHGOds20ETku+f037fBv5yf143HF0tjb4hrBiRPtR3Bg7PLOc0yMfnT3Iq6T3D
oxMoYKpXtbgKyQLkv/huIHgXowmymn5D1aeiIEnx7kqIT9STKjRisSL+WO2Z45BPOUPIn/fCFIKK
hqbzD6DlWiXoubhWUJAnYqtJaSQrdWar61cNgliqJ6N8a+Ik5J91HcxNXU+Dp47/FvwwJ8Tvz8wS
iCxf5mgPOsj8pMSJcsWnbbaZEear3v3rDvhnq9tCbIS/6TQd4WlRwFwOhS3XviX3XdprDOpQd2EO
DjsBj6LClSSpmtKYxF1aTxXJcztIj+hP6kc4tRq5UC1Nm7I491q6k3CASnOMoAzlDBiQwhCi2k0o
SnbigtVeaYkNrU491zY/+Fn+pavJiMQ5XszsRiHCv+nRjomjOMq9eodMV0590tS0LpQ/TMLn88W2
lKDL4iGO0AH+0H5GwYxXcIrzlWcVvRmeUlukb4OjwmQBb7XiWVRI0MNfIfb+fP9ALHKGFYkaP694
z2sYyab78v5l4Z5psEUTum/nygcX4ss6SNWc5LJvqivp6mQ2ysXUmtpIWCGiKoAr4iea18f/tWp1
ukulieWiv+RzE7jDOWAwNw0LZwDhZ/r/dtBot/59OMF76CCRzrJO2u3/ZNChtM163f+I1Cgi2e5y
+7rUxGaACj0XEMXENUxJlKwj0SH0xhDJBCt3tu1TwUUBgxwA0A8A8jTQNtkQaNW8yRvM0ox+yoCQ
IaCNU3zrGOTiAsRyx9ngn18/6yh/RJTIcIu+erz/AwAy8rSCqngkFzJx3AP5gJ9AgndZDEMPAeN0
hQWHI3GhrhlW8n+g7aaOWTnhoz+b8AddJEzDUmIxTi3ujBCkFNMxOf/xqsSHIDLw+XOEUMY+4s8s
+O9urmn9fOKQOIAtxBhqI6uErwIHrlkTKTzhU7r/DhlPb6l/rp+J58HY92RM0i9eN88dik3FkN5L
h2e9TJlnDLKkIchcWY/5VBu7ASVJOF9o02csUzb1sevbRkuDsyVfsIvgVVs2aU0M+NoAbgcT88Ld
txuPna1g2KEugY7BX3mncoxJgUVTKEvoH9OK/3LJmhrcx4nDlUyKRiz83N+P+Y1n23RkWyNhv0ce
qoQmAKmdjxEKHxj6nSNKeU9qPl70YlWjVp3a3IuEI4beXfLN9VRGyeptW/y9ubzb7IHuSLI9wo4x
Ky8Ui3iFDtYWyfmHi1WQuVmW7oDyw/dPrfTA7bO7mquQojoip23dqOMzIW6YzB00OVYUwpdEglmm
bMNyNXoFK4NpuriK3aqXwr2Q+VwFlv8txeczDlWuCwNsMMtimK4uyCl6iPIo/NQ3tZMCVrY4OgDV
1a55WeEk0jYzXJ7hjtKD2BatY4dMyY3nGbSxydeoHDHn30pbuPb1nwlb4RmVMhrtbiIyzhOow/Xu
qiUKt4e7OlPXiBrmLBB68wLm508sBMgPyMdubAdtRBP8KhAVT2Ka8iRwHV7XRlf35QUvKUtSLQ+D
RsGb4ddy18qFks8cbBnTV0GGMICMvDz4ECgjvn9jHCj2sS+0KbuAWqVfpsJa1hsBy/5z3Gv3ihIp
bUpCJXw/Stz7DMzl/UwQVbMs9PNf7i9kvr6SN9gmYpqOlbbfkXbKTat5cddsr626aoSAUATElUwC
gr3LiazKR3n+51TWOClgGfCg1srJbZFR+Eu9QpvDpaDZVWRELQwpUcFw0kkFvRpQc+88nClOPc3+
ER2A+CybChaROyrIRcVYQbU8yqH6N3VmsWj0tOedv92b/tYtpSb9NaZGbFNEMCIkRouRM3JnVSXJ
AV0+kHPNUCzfb8zknxxRrg9vu1NZiD1iVcRoEcbXVzWsLLm7T2t81/oLG7xTMqkLd1Ll0Twg+yux
AaCRRImg8HNEtS5b4xT5ojG/fhoK3UfbwvkwX+Gjy8XD80EoxmpuetLdE8U22j8QMySlFyppHEB7
bemAC2nF7ee2xmHJR9JFothZ1zV+5mZ/D/k2scYt2ciJKc7zDP5CnfisLT6Taf0AHRiGtj99+che
5I24HUSSZ8bqpAKm19BTogqrHMgUX8A3A+7w7XGa/2kSP7QxHBBguou84W5IKAEnA9f5Ha4c2cA7
uJ/tI3uVNOtAOajcCGliMjaP8FtLg/TAMY2gBz9BjjGAcjC7kJa8rcw/altFPzeDUcJa34jXT2n6
AAj0dkBGIV19zAwVK8T0YV871TFTFKNmp3RilhGB0UMjwSUDo6s+c0LAqf5oXwfgfNFEJKm/zy1N
xkPHyp67QquhVbDIuF442sSNppiz/FGlJySUh3HOURs6oZoUSLvitgMyl36a9JODxoAUoopgmLu9
MAiN4dmrDpMDR2qsxDJz6OwW+HQOP8r/kgS27ctHAk7CStUlVpQ4U10+kx7/vAzBtgPtxdF/Lcr4
ZJy78WVIM2PYlic262ilxRkiMt1EuSAVnsIykrygie9ZQVcVtQARa6YaehMgN0qvNHwbjrggg1EI
Cb/6YMAMqXpT5kvfG09NxhN+ZREnpbPPSxK6tddvkD87Z9scQFMKZ7YWOmxBumJ2KbAZHqMH3QIJ
2PBPlnrx3QGEZMpFI5Qmuywr5Ygsy82Rbvu/07+6cKJH6pAOQdYAW27lYpjCFJU82kYD+fyv7iQs
3PD1sJco8Phn9a5B7sTlYjY9kuOngko/9YCTIs3lwFsRr5ugPx4bvSGSER7AntT7lrmpkj3wDXek
a2B3owVP+dLjOGBBB9/GhREcxvDDMA4iTlmJbGWUPaMnAEZ1QrARxmp7tKMkGWobKS6jKPe+untV
N47vk5EmAmzfIeoq7Q9DRA83uUvGBmikYpjALjh3Hmj5UwL756YqvzwOUjsDLf9HLO136MGZZnn2
RyBAOCwlhMDtKRnyrXeQuRAXlKq2Wef1ztHxFIwQkqf8cYc2IefXQ2rfSSm9PqY5fMjfYgLMSPzA
Sn/8cOb/+G03cZIIT1mUaOVTdvzEZFRyIGJFOmG2LVMFrFm222qQN5p/jU2hRn76V+zj5l6Q+YR/
Tn2GcNELU6BsE8xhjj5+hA8skW2GmYWQ97kak2jW5Ys0xuE4Fpyho37LwoRnwwi33u6Dc7I6+Rnv
2lu62UHCSS8QR9wAuTatUnp0YyoxfsPL1c3hIUuKzHiJ6uW4XRK5AgkTn1vJS79RFPWGqjAN+WbM
lPYvzXxxaNDeO1XUfqzEwwK1dGsYaselkapX3B/0bsldFwHUbpKHXCgyYVn6r+DdUJL+6gD5QyaD
KSyHyXNu9ulsxUrJNJFj++8+tgmGsP+R+HJbeZr+zCoK4ZvDCFLUwTN7ALABkZCovKa3tyASv++x
17ebESV5wyPdkodP5psa9aTiMX9Jv4UFYRbGSqYk/YiFO9HBwfyBgzlPTV3IYftbTugV2tXJjyLa
YaaYra55f7qpk/kUrIYsEk+wSk7bc7qFzkMIQSuzgF0mnZoL391nqRi1v+nkU2ocDEo8fewgb2Ne
U5UAhlHOM1/wHMNEAasJVwDxDah53xsSYAM4LibHyDqXMMLS7Sb9vzYbCzGRB9vrHTK/vntO3lsl
VjpD0cW4vRLZlJRohOBcp2GJLk2vk7Ysfb5eh9WcBNr+X8TE90gM8/7oCkc8HUO0yx43aHtGSGQt
2y5+Tbl4NRqNFGJ3uOSn5LQLQ/iwz8klEeVebABkBaCPukNCnsRBy0Nlx5jPw9S7bOavyGbDpscN
KZnJY/Bqiv7r+N3mNwo36f+azFpPh9DT152NbeNa+0GYuWVhxYXhctHA9pFqwDmG+1ymU73+ZqN3
eW9Jvo0qjmzLx2R5YSqYwSg2PWps6baXI35RPGtGvDode1JN1rInuJe/Z7DKipIYoWVfAJr60H+0
bXdt25gDMu4JMrcA+8fTwtS4skwUpe/aPqT7cKt6Bzz/Nga7bCgHB7xSqzeejcrSzV586F0FqcjD
oOYStihwAd7BK4G7lz9/nJdNfrtem6j8gWCRn+u/fIhmOwuJuR+eRXS43qOYUB3tA1mTzJqKdsQv
GF7SVV/DG2iDy7DY6sGbDTTpaDwcQ25li3szXcu0U7bnZIdHpTHv2V84HupUxzZprMPtuUz0tRM6
kIIpJVVDPSYwhZrzHMhlDO9jE20BDgDm2W+5GT5MDbOY1wPBPg7CTRR54HSjM9A1X2Iv1znm+eKS
kJ9yxTxdrApm5nJANAFJSyMBAz3Qjg8yBHj+Ydr0W5++mXoIS+IkKLW9qbH1swwnJZ4wX6XKBGkF
kTRsHdgI8dQJRNdNkT6qkzfWkjgrYAgJ+0801jIQsZxBuAMmm69RjwJ1RIZAXEonOa0olfr4pUrI
27NPTjVg995uHTGvv6MbkRkeYsh0hed0R/vQgjcvkvrwMywGR1T4Pd6KZ33AdGKt39AqrMeRIvpr
5K1z04y0um3gN2ROVC8CVvNju/Bc7OJOE4hmw8njManePIUlOzevBoU5c03zmViajZ81Rynjywwn
wz+zEt/x729+kyNiBYxdoUOEtSl5pe75iG1YvWNo8IfrrEwyIAHpNgJW9Po+b4h23anUNrYPVx3L
sHf5idCWIgVxe71Yg478764UkRRfnRypMldunq14G4FRzZsqKo+b+4HRgTxeEO4VNJ9IPeWbkzRt
gE085wfc9lQM71kmu1heFXq8o1k4fFSV96SUMRFtkoIawR33IZQkHehga8xEGiLJ/18p+WkyRbG8
lHoZrovaI+f1v7K1us9Fx9MJJ5n3AzLJF2mZPPo/zuMayYWjtdwAVjRRu439rGiu/s3qJqTGH2gb
Sd7QCXvkTd+cebW9xD9/zq+i7ig+a90xsbMy8aB5hQgeC6lAtGo1jAcHJVHTxmsV0fob+QSzMYcR
4efVbF/SSO9yG9w9pWSgSdnDTnBAKtQYj1NygZH+PrERrewLpVzrx1yQtqLwF62szpZJ7sfg+zX3
f/0apbF/rOn8Uyvx8AKEpe/IEnSS1kD1GvlH8FZ+w4XzlWudS+aTS6iZL3Svvizk9vc+aTEMlrj7
6mueshA8IrAeMrPpoto0ojA3y+sxeNyxo/EqB8bsvtEYKqKajVoSvyKr16rLI8aAhC6JiGnH4wWq
e8z4RZex+oMnMzlipJodUiuGBRbuzEWxYVlBQHZDdG357FK5WqwgCd2z6R7azKoa4weVO9+WEzZr
L733xjUZCBtRxyZNnT4jOqceUoqm/ndM+XBUCFw8XAUBJHiFjiumU5EMSndgIX4eHDyOMzans+5m
/b5cm0gAcfUkmVAq74UR/QYuIZ9BTi/ZCuBzb8hiXfKDKET7IJrlEQHKUR1nMoBi8qSy3bc5tUtO
2UNCZmhEeRnHiJTAVW8ZNB0z1/UtninlwwRpTEBCHCD7SSkvI1RHd+axW/omd/fJ39wJYwNT+Jok
nEVGgXp6OrIgWiMjliclxLQkA1JiD0EffsJJWK6mN0bZD0z8kuVGxwcaEJyjyNPzww0atzAXNDL5
j5HLqDXlhs9D6WdQnZwcq4/uGPz9IkmwiZUcLQnj20sSIwZwl/vyGzxqaBJMVmrXhenjBuWHlDgV
vYR+sqWm1ogT3elaUAQkkgcSLQn0Dv+9k6vBzKGAkTk9zjlyw3WNAOTxWx49MNDCxt1sfpikkmBl
PPLfeckUsjyoGlcF2mweE0COr1wwHhOrCKm2b0OJNvxdLSJGttjUh5T66x0U3+6hXfdGm3KrK7EE
tqIyaDGmO9RIavkVwso8mN4DkMwxFE8N2i5shhuN/Y2BjLwE94Y38OGtqPz8QQYrTy+RxJ90hgCJ
ZGhomJ0JwP34bfaivNUEnWk1MKdWxhLX6WbISR0LqFhDqZHPh/IcinXC6zlqMdu4mS7Q4DlSBYyl
DZHZQ6GN30rX69bGNALjP6Y7dLiA9IQFsPONpj+PlLQFC2mT3oIGOEyYeLKjOuCE+GsiZAeeIRPZ
Wn09dMM/DaLw54z/BkJWc+sMHSBp2vvF9NScJaQdNtTcAEHlrtf6XeMWq91ZKzYblVOvv2OWllne
qdxUIHcQic5T5VU8WOTuV2C1K9Y+iSSeoABUE41djTSYhflEJbIYjGqNE9VFPzdTDkSCLpT09joJ
lmvpfhMt00RHmjNQH0zdIYalEVom3cZgZL91vry3YrKwCYpkqTkvcHn3rqhNznwt/f+lyRlqZKIi
Tx0X+yjIUTXdzDG1MG5k9iD9lW94thaiUFLguy3X+Qgg8X0fOz+31ffEKRad7EttjO4ZGtpOS/oX
02RonPRLAK2O4/PMS1JWlLBQmZlgA8DmVygWeb3T2bjxoI83EJSdl1+y4D7HG6XUMQVaKPn/Glo7
5cyxkFA9qRsCn3heUisuH7zRbGQZJAPUJUAKjRbrxkkpxA3AMyLcpy2yn++rsOlmVeAAWnw6OWPs
DxThwg/aNOwdFqVn7xzyL5OgJ4Z10sWxyPNi/bF1z1FSpN7ws+KlcBz5ruGvsxGfT7vpK/FAYy+k
ssGow59L3BVmYlS97NGL+ILkVgykn8uXd2XWkCpLWqkvgkq1kM3IR11pYP0I7F/woZmaOe4Lx5Lq
ZvICix2uje93D1QCZ5YVRf9VVqzh42zmAcFPJ7X2WXcBvDpNVgNZOTuYA8uBSj7aKqmYPCPxRk5e
Kfxe6+dCTF0sevDX8ti9X8W8MTij3TkmZJWF+hh7m98DClSoGAimOh8Zjv49UMxbsWvjpI8B9/vb
vcRuqflLq7vZrsb7J9jm4GHl7TJsOXBU/dv0uMzz48BC1bPhTw7c3b7ASpnLYywA68vZwxD2LmJ4
Jj8bkenOu+BbqjZSAizgnSfcVZUhTBnIqZvk/QNp6iio1kSkONP8xptpp/ogR1GflkARFbyNL7CT
gCk4azKrHgqaj50mbmlEJKrzW2EWLC10sNyUp3xGoLR+l91ajaoLUlhlVfx1548P+Ctl2WigksBj
AmfPOf2BgRvmZFMAueTrrpelAlPDBmTYv80BPXzqpmTzGTrRV/Y3gBAudEtnauXZeTMXkhzKJGsz
oyD5PKKBAQgSK3DvPuo4DHeOcWZyP1EDzLOzMgaEvLO3m3CkNUloEvwMlqurL4hDAv7MxsuM2TC9
zatDxKeuCuJCqhXoFZ6wILZMOHr2MNZEF6byI2fw1Q0thnTVqHUGp/rjBfwl3i3ry+Topf5C8yLI
4H5ksDJ0GPYhW78dmPMKbU/ww31hBxcMlbhzE3+YR0b+uzcKj+RiofeOqw8NTuCnMBS69hEvw3d5
Za9qMOv/74/O7Bb12i/WRnAQr+29BYETFfHvOLrIQJsjrSCuptBKvMfh+qlwgSMUf7c2vS+T2rQa
nXDBe/qOq7HQ5yeUM4lpIN/Vjc8joB8UmeKnRVunI92MT/X7w6GAONr/axoun1RNZBlxAb6YS5D4
sNYhe/YTVK9FujUqRQxX6Nq+o+4Ny2Qk0KeG9TV6uV6gtTtukMxJ3ujsX0Oa5hiUD8ANyuMKewwj
/Fs5jgtcMHCquWLO3087ZYcW7oP+r2TBhGSoG33af5uzgVVo7yqFrlR63IKdnEKq90wUdvcODo0s
D4LNBTVdtjvHgnk7L3upYvGqDYvHbQb5d0hjEyempYBtMJMS4BMwboViTY78S1eOFLXcm9GCVE4Z
2RSVPYA6PoMBCtwI9ul7fnoh5HlbuDc3LMdcTszCULexlX6MC86ToS8ED4sxOVBLKBOYSqVKxvMI
+XsUg28NTufaWq+A/VzmYyjGtvCadnB5FL+dULB+/aGENruJPyaeIWfm6aNi/cjxxWUsP/DSW3wZ
XKfLHRvTYLE3zfcSeoouKu4FgwKK52Peaek3PcoBsKW4/3f0vYba6Av/4CFDpdreVsyGwssbj8nW
Pze/ufFf2bE0hqVOtb7Cf54hl/AbL/xMdqII9D2aQXEwVIikGPdE96gIv1sJw2AKszBMXhexug30
/aePDsrafQRqa8W/XwzpnGrp0vFmC2H+MOCOu3JE6AQVZx21xSs1FlXehMkbkFOASsHv0eKs7XHz
L9dJ+hjoO0Nl9EUQ5D3FqBm9Did7n9ZKd6xHFue34P+9tr6VqS3NZIyYMhWey459KVH4dyt/YRpS
/+P35tRzU58VniLvzLTCmQCH8p9TdziTNRAdtyFF5mtqVdEnRn2QZZ26XuuvIrcPwiw3yHI4s/le
5S2rGpaq7KWX9gDP+aYOighdRXOxY1Faay2iw6yI3BAaqy5/F8xH+kj2bCz4gN54ixYIRNlbPuYp
nnMwOZqiuUF6iKguepAmaebfiZ9ngyf6tdSwdn9urGUJL0RalY9GYE1uttc+NWDduMjMwCDqgBge
d03bNwuqtAKy7LsMpFj4h4Jjl+/lMA+DfSs1Ux4pIVlEsFLzllrkBtvRNTGT/UiQ4Wzzf1QZhKBn
0m2Sj08cVspV4BthuNDmGORdyPVBkgkVRmg4uxVyaSgO+sbBH+hlvQ5f+4lYPReFLijjq1ohYFF1
+/KzL/l4Z7XNb26FjSYPMIjxH01VwWnqkEcA3yJOZbvLNz0ZcpcXtFFCWJRC1DST44e8bKtwhxZK
NWGpqyOprDYSaa5//7WFL5tp+fzNXsv4h8F1uevH4U68OrIooUwNnKhAirS8fB1akac9dqcTDYRP
JE9U9ZO80hb690UBmUTp3Pu0kYQxsm5NlwoUmXnfZmVRglQq0f1KL/MTO7l5QQx7z4KGgYa9s9W9
DIHfd5JqJr+dzx++SNQxR+vd9AwKNWoNNg4qbEboI0qz35Bl49e8a3WNSWnaokaoHHbmPb7RqNvK
yRIZkKRiSlRRsxGcRJJLU1ldRGbDMEefmxaSI7g7xoFnUi0ulx/EzhtvCIXYJnKGy23hvhahTzjm
0XErUcQobXQyYu5EwUFjlrkZh+rSSGuIXaEnG+0sGUDCeFCbz5lRSHOTz9P2JJSAgi0/ZFjE+gtP
a0chWNOLbXpXxOduUIWmFsnJqAacAs2iDvy38E+uhG5w4W71hkq60/Y3LxhuGgBYI8ae0u032wEk
WxF4e7S2HkYCk8F4FJj2ZGqOmTcoJmft4ZRoLAGzwxsgNzIHc+PTEVy0Hy3mSzxGTpf9gdJsVHTB
IJZ9MRRm67rMPOhQ6cT8XD9NQAcSqzYj/VmpolY3qPMqt7in6EfcdpEMw9imoieYz2F+/3v1XdKi
DATD/niCTrORxRobXAFHOlNUF4ZweqNjB9uG3Z+oWy8jfcSYM+xZ1Fe96V5RCbchzhSSqUj11LVh
CO/TYhewEP2a+DJiP4kjPBVe7y2U8twq/T4cHIzcRaeIgcWXxwWU/om1cY1SeN7B8+SgZzwJQtVg
j7tlC6M+Ra6ynyDQayZFJFgCb0lztbx3lRdVQggQj+7V+lCDGWWwNAk2ViugqkyyGsqKIxdFigqQ
/+qz7CjDXvXh5jER6DjuV1pL78kwhdr9IRm7rK3MrqGL8ghJTcBsxcDMyhI6wRa8lrGvDVmwD8RO
r2Bs1+wyx6koj6W4Hr6qYUd0KGtVxd5c4JCBV2oGqZsnTOOB9dyB3fvfP39jfOS8CTntG+EkezrL
4c4jdkjCqJc2AuS3nHxJGxnxzrbnJXIph/MW+nELUvg2XSTZH+EvAjdDBHYMSTgxZVQ+r7cx/jDg
evZSQ1cT8IEf/sYLx3TPi4FdHhtgFk38cJds5rq/rOG7Hj+dPmnLCmwgvoCOtNnznBK9pLNugSt5
Fcg2XcxUwp8/8G3/keNPlFgTDYc7/5es13PEIpz8LEycPhTRCrhZu6wlMiNRKD82YaT2kL5pRW+H
zDAFQ2jkfyFKwYGFkXsev8svkD4ph3x/10CULcOFHGgRFYHOby+EjtTcRHXo8qcGQbTWeIkfGZSI
EkH94TLazfjRL8tYUqTn5rIgy4+URxg3FAr329lawB7IaXosKpicGxS+H8ws9IEMAJ4A4XyNWUe2
LbL9kxA7sRPhAlv+CBndVqCzDv0zxJJ0XwEy7eWkMdnkCKzLFCOr0dMHvtLPDe/f+flJBE6/bAI6
mpCy6spzd57Gu3T5s0VzaBaI28vszs/JFd77XFKDCXHzQkudS4M2GVYRyxyiQ+4Wuh2u7FUcYeWQ
eiWBd6aVavAcUeiog1kMwQyYCAQQwkBxsmvFCOR1UuyppJwE8CVrtpw2UgbdFAGr1r6ErJucQ80p
c4mcghCZQRf6ef02QogB0j+TG3ycYyZbqueQKn5icxmWLg7t5tF7p0uvqKZ3ZnoG/26TJm10Qtpu
HsWulDiPW78uYl0qg9Iu3SbcN1luKAdbaMmuxhgdH2kaK8Urx1Urm6jKUTNy23FXu61LwVAIYetH
mfwMRVj35i1sX9yzxKRMiOOWpH3HRjWAtfQUU1HGcagzYD1ngYAaYBYDI02epqaTi1DGNzBZoIUY
Uz8XsFl2JWT5sEwo37GrLljBWR7Vh22bHLeBNxue9DdZU+pCvtbNp8RAYMI51u8XCsL+Q6iEt8bu
l65kwBEQVzNm3odjjIS9n7q/W1b782ptmwgKzcudOMBVFyD8+h/rgCUuvEyhJMCFx0GSAtsqTyxK
h/WsyHMsxEZygzwHvto3+BvYelljHrIPScQuJfziU+Uzqo9jm2lnBXI2Dmhfdv2vQcSMjeZXUf8V
sen9Q8T2NSS/dLmMDg5dzSkg44GOyDxBmMzCLKOHhcEnXrC2xTwW0Lvg04pT3keX7bcJp4RkaZe4
/DfOtkIU3IX2ouUWAWK0mcZgEtlLEwLq+E9Pqq/Efhb/Hiszihgu9Osf0wmzu1UWR6Fv9gsMWOP/
5NzeN+GsIhQ5lsKUQ61a7wNRFSjsjKOlAPjNMYq3vRrQPaxU8mO3eioSA161Io/AelkJIcE5A8Rx
59IZ3FPyuIOSCidLE8dZpdOPhPM4V0F7cZI+VB9HCGGByxmjkjSpvWqV5dpeMky2bC4fjH5xP6sn
N3kWfw/EaNyl5iytlA/Xh9nqjjxa9QKn7yF6P4zage8iZAX/96U5op2wVtMyJsVzt2I3WWpIwx5K
4Mkx2Rkd3J1GsIWLhmGNaOtBPLoxC/bOj3HkSZQ6Csl/cH/Cg3LHJa8k2NCkGkGOCvKKKbWfMgaT
YoD/L+wlEgirN/fkHHZUqZKrrIA58+/eFdrM+VBWYKdWP1PUetvvT9ljsw6EPdcvqS68JEjcV0w+
4INEhJVySsIvoOg/fGwE/vUwM3nRB/98jINGa1oQG+3KZJdB8jX5bBEBXj+p63o0jFXvcx8cLKZW
t56B/jJK6RV3wQQ3sDR8ilX7FfRcvIbYKlRwOR6MkStAldBNCSLfPlYIOF6omAxul4b1n/jW8arq
0OaBdxNRkF8xc3CQt6zDKZb063JGB8RdAryCbUx1nRYHa5sx3NDVu0CXL27piA3f3T63Lxr4ncW0
0YOuE254RsFepl4D/0H04PSaWJ5Kw7uuPDCyF1h4CBQ48xpYl2Ttfj65EcZ2R+DqKJFfScGA9Dny
ducvVx66349GzVS37E5oJbdXNkmhoVkVRT6iVBUnxAMaosS5LdlKnwjAcFoS0aFD3JAlvUSVGX1X
wiA6I+ylHLlhVCKBAL+9ccPEgqzU3JZqx77GTtUL7DAQWyDAcP0f08tsHGm0/o6Rshm3340+Zu3i
yVWR4I0/s7gaVOjAk91NEtxXD8G59dhxlxcPBtDeupOONyGyc0LtoL+0fZ9VOZjNIgYwk7bWBexG
/NGyNgdPcHj7MnncnsqdcrqziSxu7RaMsfDHNQpFWv5VdCEcRW95u8jNiGq/5Q9MFQsAvuAP0KR4
j/8dx+mDUaDrcsYuJ2mtBsKI6Anbz5tahfYTDkAtkvuKuV+eEzpgbU0w9P+X+C8WSdUhDmtw1GAu
aGReRGWvhxtVSsR7wIOjRk/uf/xe2fD9t1j31XlQdFVBnNKPJ6R7Ea0t2O9cF7vx7hbNcvO7Apk7
m3SWTTSwgFSgRFqQVXCkBrrmAGlke8JzdiHwTCXzHWk4/ABQUhhuKSZXlodEyS3Ovkwb4vsuXIo1
B6QOAEkJPZjAzsGsGdsQbE6Il+dr5f8gEmJ08t2SGlSrwj1I+PyI1GmC0wuNGZMjbusTR4xo2CKJ
I3KfhEGb+vUM1hW01X86KmZ3s8x72S5Oe5b68ziaMSxvdqHL3uct5DgZju2FJenaSnmZPrc3z9LD
impyJ16Y3rObKBie6P1kjx4gnfRHNcEShmKdPMfi8PTEiiNCKgeUzk6B8ZI8j5EjZOZwF99fIfuO
zsKpI6QXyiwBjw5/A89x786GZVBAT/m6fim/V3Lsr74rjXaRfsTril/BmVM/pSDqTzEFvqCLVj/Z
SQN8UY9Tb6FAawl4MyUlKParVpp/HIWibIxOZ+05O5PwHyJ7VN7Dr83ETUctdOwCixQpuEsE4wEU
GyWBtA6yqsc3U7KMqPODoEl1NLSPfOqV6Xra71JxRkIBNoEycGvoK5fyErKFADkSfbJwVOWeGevh
oJKxFqEtQKnvLmr/ZIrceZ3JIFSVfG+iTPV5oNTKumYjvWBRHCVRzVTpwx/5pbYznTrGWSlksEKk
hfErBVWaSnTsR9GHk+JYCnzGxQMmB0K0r00fH/vm2YpVG2S6QNIGEeaHb2YSGsjfkA7Id3XM8Qzw
LJrRQ8ubkJvN/iewH2RC2fA5ST7Gqg7L55cX0Ns+5e4GTYiBadDwTYU+oq5HT3lWSYj/re7Pugnu
sds41XfkMmQ8KU8unLUdTkgYAwTAPvsPMTIk0cCDv5+WqrmcLIoe05NipX4q//ZjPyB6XX/yvmBb
9qZb2R7sbGbgJELJWMXI2g7c4buLc+EN4CAh/qs7HNc3SmwVmfJOPHg6UJzmXUAIPoCoYnTnK3JD
DUQdj+z4qSff8aXc/XuYPjmuW6fboY1nXPLdte1oyA98kiD1nDYji6E06mxUc3Sg0j6hUQVjn2r5
cjMoq7kLtwGpdqybEeHThsmqbXtXVI9o/hV1jk46vBTeTSno3Kf/iCtAbidAa23hu5yLJ+fzxAU8
FxRfUp6mUMHbYGhLPrFEs1NkbSR1hy8vI6dN1m2zk/O2BzIDgcFkdGrFn6qQn2pNFTR/u1ntfHwl
2IclUB1UhXS5QIepXdFz/HRUouOX8yDjkLd2aZwfj3+g2BoGnBUtP7ijRMHhapGjEMGpW0yoXHhz
T8LXvy0SpuWWBoYSkXQ699F440YdZaWx92E4BVBNpfEPvB9bxVGrAhG1rCy5kYh2eOZRDxhOvCwK
ZkAeR2xdmZKQIk0SIC1CDM3vbdUuPQ1Z8/9xc8oDpSTYM+gDEOs9sD8OyV0MNrcFtjcedkwX5CfG
hbDb46HMwESmFMTIn0zfqLOydenaN90vlswhKoBPsRDdVTDebLWUpuTSPG9lcTc7jPDbhPmxfip7
Kye8Abx/Ji/YcgtLLPXxfUOIVKtG3eHpJdn5CkmkzjbNfCm2QG9DKcoBBkBjN8Erixwkv/RhUonM
Z8t3tLhlOMJvYArFL/9UCv+MmWzsqDnLfqDXAzAs1Qe9SK4UR3WZRKzJ1wEuy/XrRF7Of5957KYW
Wsi3sFp0fHkS1As/oAKu8J3FIvOUrbJlYTPlM0SHArxIZvMuTu3kD2q9aJ5+mM+D+m0wWvigZyHt
iD71M5yBFLKX3GWT7FYquT4q3knFSWR6mS1/1/jsLHNt7cP7F8AmbNeAsHcnE/DY1acmZ/VEdj6k
3b3ACEXqlMZ3tf56ArqoL5dIGvIBvvzejn1Zma4LmEj58j5AS8RCQjvDfSEF5K/y6Q/0FF8gSfNn
OyDkokJIO/F74hR/O6hRbVVGKeJe7aZmb/qCNSajnHgX8j1WocuHXoWNUNgXSbe71hLB7WnFEPYy
i559mFbe15FM2kdZpF5M0GgC8QnkiDWnK+EIwSHw6KvzBisrJyxVmcRwv5CC6LpG1uyiz9QK1UQQ
a+WVmWMc9VYrMapzl63b/VzJU9bh+BZuIMrmFrCNLiRJwtZK3CGavd5jc/XZlvDIa1JfEZIUZGYN
AIvvvkAJKFnUtkH4E9iEl2wK+KylwWlwfMJrONx2faUYql4CKQ8tdW2jWEpC259H6GVmH9XEyAB2
oWaVS5rVmw9Tlbh1844CgROaL5pboivmj011TZEpVWqX2WoS+8Ok92BD4C3860Pu5lbl4evYkqqO
jLWSuC8hx/6CQYsgMxZBgvgn5TQeeDsTBDdKmt8US/Cb3dtQEWoIC3e1Tx2exu+0F2Ey9M6rxY8g
PLq0YpO8bKBzsnEmk1KrNBqOQaUEL478xGssbMCbUxG0X934UXA9cCetFMX2HQ99wmG9ohOtdSC1
U5Ji48VpSL3yO4diKu7jYFirdH9BATpwsNgaYJNdU2p4mr2WND56tyhhXrH3o7sd39iMRcxRUkDl
4k18uBfyhdLS17jgwZeZenOKrmvh4FJsV1cHAb4qYQHR0qmLLKCUMClxwXVcl8ctB7IDlJ71Ae1o
ESazKSjNES7DKVkV9gZN6/XXC+VE7nH25hoP5vX9gGY/aUDn9aoWNVVNls4kS5c2Kvp9pIrrZxND
D6ppE77c6a/rmUnHoKNo3jvNiTf5xZO4u7MbWp4yV1O97b7vtEACOAWxP0fwsHvZ5f+Rd0BGkwFy
IW5EtgCyoZT8DgiNMHG6ZMT5fbWVwd9DOxEunrBiMbP0rHfkPCAgwHBhUrV9M3fB9CHcFOK382qM
mYS3GPuHn1Mx0/K0PutJdVTdbv8oozPUmbvF6T9yAeRa2wIEqzcpCRJFX/DG80shpPj52Jziub3/
XDyONjgoWMtaV/MHvrSdkixjAlXoOU4ke7ybtkkWQz7Gk604i6kKf8tsPoPm3lApnJL+mLh3K8UK
rcLrOrBwbLFrFV66v9rNvPYu05t1bYwPTwxr5biI/Eif1M1eyN690D0Jop3B7hlIqnU0k4kUAdxQ
MJf7xPoowG9/qIQcnAF4L39QDzRjl3J9kke+w1onxS9Za/YnyMf3ncQaWwauwLuNXAAZZUYfIHoN
Z60CjGhc3SUIYUQwvn4b4Ktc0tLs6tBpQHsT5pcifUFtqBPdHMsYU7utXOFTO60sza/eloFXOVbG
JLLQnLXLwAiiOI4FrPG1oLn3bqJTPRuHAo113+3eogowyk4ly/7znL7XOaHGw9/cVKicQwqdGoyl
cFFNwMfozG7T9hYcgDFuGpudZXQY7xb/yzYxgoN+FdV19Zss4AqYbJnrrqdR+VipImOKetIvTccc
BiE0xiO4cDIf+33a8getWzsZ8cob0ZIvOATdA5SdFf+FyDrnKOA0oPT5nU2A/b+qhD3+kY3jkTZB
jgZpotTGUsJK7iFW/J0xrE/9Qsc9DdvM/Muw4+84QwdJf42AXFDrYdZwU0a/b1R9tKnyCZwELcJU
Wi813orD76g8tPHIcOnACxpUm3JaLbS0DklWTxqhSSWKAC0Tu+yT7WkGyBLXH4qsg8CKUpOwUaft
AERq7XLdmVO5axa+Yh7GqqX/U/xbZQ6CpObKbRCDZ1qcIRiKjjWcbmFquaeyhU8SDyeNwl4RQ9mK
OoG0kLQlB+SreK9dAPt5nxB4ljlHVHmNXhpB8wp/cXcFlUSnxQ7f3H1i6b+VljrqO3siA/G+Xfdf
Qik8G5OFJAa6w5B1V5vANZJlkDW2h7L0CxFDeMpQE7H0LHcRe1Mb6KW/JXf+kKxfN4RDhL7JPWCl
E69N5j99p7jR/GAaHVbUYb6U4Z4DnHtwW/6+q8pIN4xWNo5nquQibBBi3JfsyDfFvqcLqXmo9IFO
Pp7ckeIyOypohqJ1RMJHzVyF6poI2InVrYraHE6D1W+MuaUyH7j61TAlOA0eWWD/zPmorshhT/R3
ydkzuFkzaAHZ7MulV0DJkP8SBvquMq7ZVjLDJDK1U4VmmMaQf5HX75clm+W71i48G61jUUFK1LgS
C9BptjHhchoTTlF2O3zd1wKQHSEr6Mjp4gkwyBOaNK1ErNQECPdJt/pzKTd43k6Jm2o8vmzktgnU
RA3B64cxrj8tSK1eLJVVgpmVuYpckLD01Qet8PTG/3x7fnM3yp79J9icZ3F9VSpYPW12mv2uBZ10
LLIp1NoK4qQKiwcbS1/a8VZRRz6tkjCrrfVf9LfPrg/8b7jO2kyMQGlCh3r5BXDQiLRU6YSirDra
7VCyCaHVN2oBuqlBg7k4pDvFC7dNius7C4a7gD/3/M3zOw9sn/rRlRthz1d5Srqig31L5H9E88xm
ywkosbId5bs4NTi54vbcJSuC26yiJOwjCQhGEOAP3wal7l1He/Rh0AO5Q8ia1TN0aG+SDSbOX9Ol
Ba/V9gwlUT+x6GZZCYt6rVSrp/QWdz0wIgcnccLmqrSqYENtI0RMHLpVimazTgWj/ptK7KQoQxuS
+47CiXqPg4K5HDLlDho+dASuSYMtf00esars9a2+cEu5fP7uGSbWE3kPvF0ee9KrjHPQ7LoVKm0D
JsoY9Ft0/LV2baOYNoAmcDmaf3v7bKkZReIBbud+wiUYdMyv9DN28wdY02JavXfMYt2D3JK6zyNI
5B1Z21qav71Gzo4Pamvh1XFNPmEUYll0tl7Wyp7SNJhLWc9leC3Dz5gmUfqEbML7bXaG2CNQiNqi
OLRVtzfWnH+VAWKZoSxsRUUUo0Dsjz7MAUJP0bIDzWKOmQ7NfD1hSrh4oaoR1OUWB6gjzIDZFGG3
tIeLLrcM/rI3uDGmIo1mC/jIoaj/548rAD6m5vToB2O0xDCmwl7VhWl1IwKH0FRIBQz3oIkXN/u6
rJ9289xM/XUV+nCxcgi7tEzI3baEVZt97UHAIWLvmwHaRiMZfVIoqDo6zFq3lYsMtoJ/+C5rSLU5
xZb02bj5nv9iqHgyiqf2nYVXxR2njP0PAMkg+7oVddCqpHGJ/Iui2k0JoyAlSeU5AV6CS4BjHg17
lD3a+z4FuGqmf0W/rf2N9esl5SdOZjTPtVYceaQPBTaL6qjwM/GoNgY7orfevlY2t61y/KjkbdrE
W3m9ZtokqHrQgYrgMhDVNqZfbuTm8K8w7LAIcxCl1vIExJEvsyp1wXZJ3VCR9p/YBgYaHgiA5ZAe
jdtE5NXvyjYOX3c+I4Nt2l88JrEJStaeRFjimpuvgj2yL1lSJ4Rr5GJ+uilDK15R1b9nsSuWzsE1
Pe9/Sl58lfah52P+KnlOl+30+nEQPinf0pe0e113LyysS4u1q3bA09cCxo4I+AgMbRNhNOcnvxKr
HR/pfvSGkiAKqnY9PiNQiZ3ZZ4MsDFMAXRMS5s2BIDaG/B907CXksM358MQ0BWIWzeKR3e7+dAt5
YVKnV1EJalOpgRwoDokrT8r8QbybMAd/9y9ywbceEflWjJJJVncrZxmdwE6Cbipkui1uL9RDDqKj
vsRS/51Fz/o9CGxQXsou0Wncuye/oiExtw3/udBpSe8ig3I7XYC6q4UMjhyI4tkUb+kVVXQpcqeA
T0Jb1kaDox9wyehuPCuOcu6lKRgUPjwNgYpCCxDuAw/4sI9kg63i49KclnJ0egB7/e0/1Pj16XKT
fdw7Ys8ng9LzXfwWg0TtkziAc3b6QZ6vSi9OnlKAWYnVUj11BKr9KVKdB9lN4R5oYAL+KECS+IPP
bt+ejOeFGEyA0SDfTBL3XcBV6gPhUclHxMVrl94BeMRnQYl0sz7QPxuukCPHNtT3b2vTonORAM9j
5LN6FMbDN3EnFJOOv9gci97pMqV0AsE0b5J8cEk3weC0Yq/bU8T0q1u4wgVrkElG0B+4bnbY4QYy
JzJmqMD+nDzxKVPztJIwGaADx4ooJhDB1K7SVu/ZkpU7YsHNvtLQAjd59JR/6+SWpjPiTJjwYgJY
CLcmdvKvTDttyp6xvSTlQXXiLBqr3ZceK5wJB7FjdbJ06Yuk4xsFOimlioqTN+0JmpN/9eC54Tkk
dc+FIMCRUygDW8LMlw5qpvTP2+FqcgfkWkNtVRfVmPzKi3tG2dzSr1iP9YDLIypX+fOR5ihW6OUX
20sMelVJgfpQ//N4FEN2KZvQu9XAb8JceaEB5eHwu3iNM17MDrE0KKG8r0+nidEzj30e93sTJg/k
8DWiXsbpaJbDRAjl8Pswx7oIDIu7WdUluAy+PR7Nyn0acW9hi6gWHvwDVAWR2eMC/oTPD68QV2sS
CSrMNY3ZvsXCSRdylqtIFjLUGRYmsxEfZqpuA1cwLmFaMxOG5jU0NOYq2X8i3BulazinT38O7mJ1
bY5mke2p8Yndifd2v8E60r9f5xLEO2kVe3VV5cbvz1MTVc+cGmcPLPmIkBucOwTipWKXd/3pn1aR
R5R3BIK3oX6RDAGdiDV7HcbH34DMf/K8Co3Dp+JYioE6nKPhBaQ7ye4uqu7/eTPSGKU/oQnj7FrW
NkxsPoQHE1y72xdqAG413lWs+KmcntspgRlGLchO6N2LTgzuYUZsV0mDiSV+n4e/NcLKAyeDbblR
WWP9ePI7zjWkJbQXajk2eihzg04Rs16SkL3faQjor7M4aJHFMhRAiUtVKvvMzFudwD+n0LNTyc1x
fMrHbeui2rmtdmq43cIyUo6zewQ3rpFcprqXGJGjqvl72MsSQTHILalW4pxTK7FM+xQTC3H19J5l
NsspPD3DWdLPY22XDDEgJl3MiiArrDwHyqL8Dse98RgFMsVKTc+fIxdUrLFmdlt2cl5r77l9GrcY
ack/kyTy6Rbl91NkwFtMeg3OLsNDsOVIsHzt8cK3mDCLaXOnp9RMJJU9pUj+vgK6H49uuiKBz0bP
LnWUEgcWENkS/96yPiC9UXwA4tULpfSmFFzPT9ZjcYVDFX7bHHAlZ9yl66pP/VmYBwYIRF8/Tdsf
5uXDkHzYkw1qCs0vC7dMgSAxuSY4FbKqxNNfS8VcmMVqV4Lk6/WnSlVORp+uIVnFlMqqrDtT7khC
KPyaXTC8IdgQK0TVhQBM68ujylY6cIGkTtDSeOBhnQeLtd/rNcC1+/vRzw9+YLdv4lerz0z6TGUh
a6W67X3bB58YGfrAMTEmaqnMC8fIge/bA9jKC0j2CyL+FYAvxdPQIPTZkFyGRVa1h+clONadAAJl
hvLksHpZTwpRKAh50GgjvRvx3CqYgrPYhy61Q44w/MHspJ2dO3Zy2L7lgZbi5Ssa0mcYwGjKDAAT
IGgRt8E+4jfL0V4INLGSg0S/8kB9yw6arxOR2EJxORRIUk6EFy6WNGesH1qdKfvJ8FP330VwBFMD
n2t8+df1xnK/CUgcz2QAe0TLN4wQiqIgf8p+amgmH02DJYBU6WBVQNpEH8SjMzDzJrMZyiNWCq7D
UuFMJG3cck6M96plxZxISwKhPqM6re8RxnV1qJlXuxxDOT/D9/Jn2CSvWTvQ98MoJtCMpEUGqYD9
HRLyDrxf3SCKTe0lqcwSnl5sJnKkTfmR4Uj92K/DkLa32Xc76U88owmOKumbKRjW/kZBAjqzrD1/
28BS2M1n1t3+Ztf3BjpR0vRcJU6USvvIaPRokkEzgh04/2ybw0U5cHGksD/ATpenXHIJGoMqDcHg
m5BFJeTkhYtNqr2sbpqjTvrZtH6cpT3NedFP63fXWsBCSKTqPI4zOz7/cFtwE1clNqjk1AYKlnTi
+JrprDr4IpVtzw5Ksi88z0KPdrjvvTewBvlvcOtaqDgyLLqilZqKMrHO8gUIrzOOiGnzjL9A/Hdi
ZGY6QM5UaYN9TPCoR0aO5RTt03lam2vjpsFQtoFHyCYRyxibGVgP/HdQr7774wXYbOyQ+Z2rUaEd
D+5KmHC2n1H4GPgTIqtA3Q1JlEKISVNMUPZ2pWw5TnSsPqCQM+ZDuanfrD3rl2lTSrwBKbuc+KkE
mOwrFp47Lk7lgmK/r3CRz59wodAgOUvg8iFqmvGqftfcDkqY5fCCwBw+Rdhs78N3+I2DPoqcOV5v
61eUuDe2NlYMQ5x7Wgc2N92Lp/quDKhaqX10ki/6SxNiNeZTvDBC/6MgEE+uzVnUdbt2Sx+knBet
nyMjSB4moRYRhZoVhUEv4EzzNRnCekVFeJszTCrNMYpJLCbmQKZKgViYbVURdgnJxkivhxScBDgJ
gwJHS9OUJSJkDFNkw2jFn+gW8+DdB/UwZjzvjVoKZzHGXW0K88XZqDDPt0SQ36x5Q3Y5k5SvAcPb
2DGV64fuOJyDibcoi3btZBMWGjK4pyf2jh64lJNHB4poDXZbGrxThV0kNWm6bmgxpAoPw+r2M0WM
mUPC4Kn+80NB04x9Gfs2Z4Rs0qkKk1smc0pIB8WTin1kYU3AKdPh3UwxGuDRNyHcWkLu3qCDTd9Y
rShI/Rm6F2GXTsxuOVd76708imM6sDPEj0BT3xa38+T2G1yWGBXB7BjYBKlDlNjX2fCmqdGj9UIP
86fWjT2Gkq0NsgHhAxkV9v1Dz0huJybyUpjZZhWjxuWgJ9TVriCme73CeRstVAwVNYzjCZ3JPaqb
BodNM2NIhbN4HXG0X6UeI8rRc99rbfDY/9m2fn3hu4KXll55+GZE8KzVIDSC4kiWVNuklbMaAxwe
pAYxB0BidkQCTm39XkNAqUAyLMWqHLxN9ks6ARjRw9eCDSKRB8aQ4Da2coVz9qn1dWkjOebklYuX
7rso6xa7V7ZlYGaPvl6ehXy1WnceRhjJEKpjba3lzO1MYtPSXnuCeC7wn2LXCeFsN/6bAxq+Lfyt
EVwtrVlY15kw2al3XehUAFxckL+J3LrHS7M3xCKMvkfzAOdphqsJ3Z4F0i7oc1ZgogasOdclHfsz
uUkf2Kfi1ehVOjl3gpU+DZZVODBHJQ4tRE7cd/3LrrTraJe4pBsdhSgakY46+MBxcp0zx4wRZAY3
6hc47I6V35gTpJhtO53HQ7fSJAEAK29fMyz9XrdOP64pNOUqTbdRsyI0RytRDSQ0pG33QqDWFSPe
c5zhQBP4tkkth83ner2czfQ6YwAEzmSkGWbXOqQciAgZCeHg5fCHN4rJcpCoh54vVPlaSAEtqcGV
qATQeMcYn6A6Hhqn2DGGkkHerUwl6S/zGU1kfelmtW8Bu0qrfWypN5QIx85YBbE4IfzfB5bJCCdA
zjamzN0SvBsevxXYJ8lghMn473khfqd6jYnHugHl9FsBK9i1Kj6Ne9xQj/nRtYK5kJ5CAKOedLjO
APHSKaFpDzMBrEo4ipJJFHcy49vZ8R/mztt7Fpnd5rLgmRYe5aJwVILsZLL0uTylg7IOxiUPmWIX
k0C4NzapyxFjp8YnUGGZAMss/FRBGGrhV7GmbK3NYMRNu2KcH3XhVRIF8/0+olE9+Oal94GWC4L3
FedR27xx+l4eOd7A/QgjC24HfeD2DGIGBBt7TZK4jjoeMqeMws43QBXqM/VlY9d0Wtkksb4Ue3IE
aSz1Lm0LTMoqCDLD8b8KrYIhkhqlfAj6+98QnyWHFGAlUvNj5zIgzH7q3Cs6aiOFiK0DPArWtlCb
m48U1XazwxLeULkfqxrw/W2p6SxsqqE8dN91EIRNeWSdX8uX6GWk1AZbrEH6MbvgoN2INeAv1AkS
hPfbu8jro6iYXDyUMiZ65rWreE0D+9IVLxM1bYuuetSmWZJO2k7YkA+wcx2QhBM+nH59upZZefED
YIQhUb1N597+09eoZHAS5E0Nd8QV9Ktpzb2Jt4xcPogv+lZN2w5M0QqKEVW6EIfHtuXEVjynxhbL
Iy7TXnZALIs7Yts9J+O8SW23++LH56g+ju0MKHbLDiEN+qI8gBqO4A1jpmN5bDafNZXkjd4xU3Ss
bVLlZvZVMUWpycdd5PQ4XiG94deGo87YHzf4u1pZXJFX1zRbJ1365iJEL1p17gRTVuRIbqZl6wD6
v5d3FSmcRavWe62iHZMbqLNJnZDfnquS0nkrb+qKn2TgqeIOXQqQjyEHd/2v2m0qN37dTaVFh1JK
XxU35Dsdc9h+urHGNvRIOmM/uFzHP6kq6eQU/oxzyXlN5tExDjv6/CjN+S14oWzyfH2hw4/rCoAl
FsRnDedj+KYppjPO2t+gS9EQz/mm3UrlcfLZ+JsjnFQHOJoXi31Nuxx+SIvVWNR/tySG4aEGQNO4
tZBpGi4mwAuIoFH9NTcFWZOPMce/mMaiYsc5UcHTaWQSx+1FigzPF5rpMebYPhh2qy8uRkXMBwcd
IEhpi5iPsoxp3CoeThMBfgdHQPDwTMpsLOrUtVkPja/FCOvvmeyOeQxa88fQ+N9bzF+2nYfrjmQP
dzZ9c8fvXj2OZwK91hv/u8lYXOqvrlMdgPS6EyhwzciRL/uKt1dBC7GOoEN8jrXhJ3k1WtsvlYAO
Lx50TjqfG+fEFEOkbv9YeYSHnalavDDlxnyDHi9YaGvl1RIMJlNUDqpxASAAZ4q9zpY5458Q6Ueg
irbJQovweD6iDAdEOwFamppItpLbU7tV0aeHIKmHgrD4xrk8cHXeoTcj42R+ajWs33FuewtQrlJR
b/43IhZQJQCP0JwpJgMyA0o0IEXOPu03AfmN6Jx1dozLuTFnuELX9w2QvRW8tDjCdr+gJERMI+LR
4QsuOR6CTqzpyRDZvQcdwbTLZLLO4hcU9kaPqGl0el4RZiayYnG+WdddvGQvwRcz+3KAQD0xWekk
c7JIOhCCjNH1Gq+f+AjBCRk2HlxX5u1r5pcyIuwAQzEJh48Vgcj2jAQbxX13IIIItigB1IuU8mNM
EkcObIfSmc88SOXn8nQf7znHQeLQHvCZpgBEcF3fUR84ByyNNoXgC3OiaOjhVC4ZS3dfys/RGbeZ
AZ2oPuZ81Krba0wQBFJDy7ZbIcFfQcnoC7MuZckdCGWtJMVXNxkBgBI5VIS/AkHTjbfS87WCJQXQ
jL8XBX/iERwtKo+JfAOP+X7DSfCjg0E0m05cMtx5beDkKjV5Uutk8zRx2o+lX1E6RJqV6P+2qxxU
dZ52KPkk9DKgWzWpOP4ERSp28GGCuPBGf5zasaoaLAuLvJoaW1j7ok34pn3kujBhQSKIIED/IR6q
F3PKV6wAWnBc3jDVhDGU2cGOGxtE+QM2TO7qXgBUkG7e5kFNOYCtqrgZEMMRy++6jiGQVQxNKIEN
ZOHhnqW3YO+QtELGUC87fWBn7gucAXebK8uXNaTIEPPKjgWJeF6qvbYJQ/i+XrVVh0wt/kaLYa3K
ZwW193085ktH4XGVXvipIa+7OGoTkWLJIRqM1qHNFJFJ2bMeOOrwmQFtlqUPQR4kuEKW1M+aE4sU
hfORaF8eiEeEPEPtF2dL2X5VqRITutv+ScHaK7dBHgowkYLsPjytxEt17ha6t23dYEPqpeCiYMWa
w49roYiSrkPLZaPJW1qz/0KOEGdxNIbQxmjyEP1LakqHFxr7X+E3/YzGKBx5S0w2n5mf4HzxBH5D
4ufKDUCzb8BU2p7FPW9D5HycV/jVHHGO0YBhUp/uUOTl1lQiMRflQo/B/nLr/fl8KkIJgcBq34Cj
pQH4KS5ME/fmhbmjDSeGdN3KsDqddorLuvCwhRjjbMyNbUlNizMq1vio83BWFWg0OIgLV2nlze+v
eIeGtmlnAddVbMuYl+UTESWTbpzayw63MqF6WPO/al5obYGVDArGn97f0f3PNavFH/dH1xd47EvX
56RHKiuJBcIO0yCZV5/CbT9A4gsWsMq6NqnfFMeJhuDxnoJb8tbrhacrHGamApbCyGKBewvItkNb
OCQesmgUbym9OyrtWIeNDeYyUC/0GeAjPC66XpNrHUY9L7QyqLDC08athGUwzOHT0GA38ezrpvCc
yID75jVRdyo+1v630a9cETzBpBw4fq7LMtEhJVz96kWZ99AOAIOY2S4AzM7c8eLC1kJkyykDCXh5
vweCpWEo/B00Jd+ZsxJkr71alh9pBujgfpcJUjPlb06zNhYmToUJO6XbUqVcFOcXaCITHPCEnuuc
WMlpicKaGJVxcfRvTZOcoWlzxvurPcRLWyyAsdx2NMeoLEBadQuXAW0T7ZQNjFyeZkRhF8SHKeG6
bJ/gwcViL58QHXLOfQb6itN1IO1PY4h21EG/WftLRHKIfsnCBMIB/Lja1XsmEoOx7hpiwKzloGfo
/nlBrVTrchpl0JCpyURa24LsxiJPgI6MJvIFos9nTn8Xk/dYfiaFXW1ubAMRLZjr9o6NANH6dMX8
oZhgeiJlJ6tStQtRgf6GlWeWqzaTBjVxg7EiULcyAQOH0Jj3tsPd+sfRx+Fx7gx0FfDTvS3aV3Ky
uOmsGouPcPhR9tene2yRNW/WOUbtw59MA4PLr+y1ld1Yczcfk3xiKzqgs1uNQV0Ki5TV9QUq11iK
QpK8qb15OlSKN7NguIN866opbGBxpAJznCzV4TeYqdzYLkGDjcv6C5il44KCzP3wUfeWLkPfhjpB
8Zf7VasSY6tR4I3hgfjoBjF/jmf9O/pAMGVX8UQ8XpwgODdP1zaALompgmMvw0VAp+rEI0J7R+/l
wM63N4Sk546con3IQ/QxlV1bcoTX2W/Tzneq/SGSlNoUF6dua5Y2GZ0DMlWuQOjVTjf6mZ6QubXJ
97TUD+8oOUbwwAWEQwRVxXlFJQMF06WghFVQ7RuPCZWypcR+VfdIPiJeA2+D5lTsRe1uPwTtCmPK
bOQixjgiIcT5bbxH8W5K1AmLp1eKZ7ydarj0VUdzaPuZtZUTwom46VGIrEkNVzwA7SJhBfWVMjPz
qI9yLRVEPczu0g2PzQ5BVhrx5VdGhxYs3ZnraV3chW+fgRgI/BIgJZpHan6k8yp3UUF6iwXCfzts
WwbHhZnYh5b5VoAI01q9tYtMKwmeS+2EaakUYXfCEbaQ/uQCpD3G8++6NWI4IDf5NSvRYfpyRpth
yzhO/4d6O1JkE6WKV6GawkvQCfxFRdHtqNbu4eEEIR5++4fbtH10P2WhCjmXTKXzobWdJw61eQLQ
vAyPgWrYiHP7xGD7FWd89rK9rBgZ7WFvbtyYz14F6pb5B71AL1GW1X//TR3NwM2MSBLJVBAkeE/x
xxANZh2a6JTzm+7NP1oxxRyJ5Aycx2vaS1spT8CJwvJUPVRETc/H52jiyd3PenNIFrh2wdmUX9/I
NeiRvkQYEXU1zxbd1bSQXXlmdS0nPiQ8YxjjUfeztku0BPt3om/dN9tA1L3ykrrdHh4Fjyx33ghr
UH7WKST89skDZditLGlndtRzjI2TdrIRGMtLdPTfDSJDiv/a/5r3q0+CGLqNuLCPjzK13lCoypQs
z/lTWjZGNb/+CRM3XA7j8G8l7wOYNYP3cINcMF7MeH0azcQHrgHmZU1izHhq3cFojrDUFREPp+2b
zX1Ze9AyxepmzbijIhGkRYOObIojWivbBy8a1aLDro3ugs0GqR4fMdfWr6sZmxH7fKX5GqAMDG1u
D1vTQyyGcLlEkFE4c5EMIfQxwu+/xl584A13xxgOlVune3qbcFE1DabG3ocGmZ/6x3irkq4vIT9s
tzKJS1UQ3TdzYrNAfSLqrnMZVuUH9YdNiV5KoZSw3B7TzQ4HewHq5qxgx7/WRLUbF00XR4fbjePq
zXIQ2vRQAsEUPFLHnJNrU/dvk++eeCIXM/rqGhWFKPa+kVJTY1Pp8Zn3D35qbfpen1zn9roq7Krs
5RAAR2HFSwe3M/QkY9RqpE6f2XDBGA/fP8qkMqSSn7o/JQfXBTcwOoNQNn6upCnjJOh6u9DvvBZN
FIYQ+hPB9sz/AA7k59q81tz1zHv/Pwtgw+ZyHKqayCptlAeX133kEIQQ5LCBSr1Lkc4yf74HhFwz
5OAZsySiDj1YP5CCVdgUVclg05QQjThX15/D/AkebBOBAi4GrYaQ45dH4NnFpsgW9j0ZA43AlwNI
QeEfqEzo7IgBy+XLEQiY7wlQGG0E+lGNo858NLq/wqebwL+PyfdMGf3bep6jyYY7ngDQuGhCoOjC
Jpw/cUxSwRkHzLXcW1Rpp1KKtVabWphPhk7DZIUBCKdrZu+KEd5bnfmzZi6v8i92+y9lVK2fo/I/
z2fkXGmZqAEREG62Y0ssMqXnGdm2VET1/64G+oFHX9kdJ529oNJETymwAVwUy2ORUtjRtyH1R3h/
sM20buJImgFl9Gt+tWPU8KT6hqK/h7N2gMf66tBmIzrVNOuw8P0L77UbKEFSsyH20oYs08bszLuJ
+UqlhRHcu0xV1scTTYigOxTjKeUb+bJzWWC6/qorHSk5nqjRkrLYpU8XKgjghSlVBZZ/pgHogGD5
j8yhEbfkykjwOrqyndeC73Jd+ze5XKsbtvralSLlEHX3gSmCyBWnVVUuHAN8SFuhp5mePtmkBEBR
kw0nbrShPFYKFgQatQrQwxWB9NfxjBKe1KEOUGbKK7rJN2d+dJaCQ5Rz9crRRnTx+XbbTOlTx5cw
8EhMVwHBgbN3sK0YnXnWwfY7hqd3nKvvZ84kvuBLXlt4KebP93mUMvj6YG4swr88+oKrwllXw8cJ
eH7LwPY8AIVJkaTZ8HCQg7r2qI4M7b0o4DcQrdwOC3uevphyrSCMU9e6+nrlw93guHQPr2pzE4UO
+EV6eCYOKNp5sqq17YDX4EDAkCOXRS5vBimRLtObXAcQjFfSt1YU91rO1R5vWywQ3E7yB/LP4B2o
OkHUi2x908XtKjTXZO5Va2TBkh6io1HWPwel3nMLlfU0YBGg1yHB0bSyrpn5lMGzkUVfLrPUiSHv
b+xsPHB4ziXlg7pBmD4MPZ3ZH5bx7lXaXWnOcm+qWXOzeUcty4qFJ4oD30FgAR2KfPpVx50MLxHl
h4wGV+S40LFkLLpY7pBrccxK7bqtaa4W2oJJIZmGAeRWy8qLOr4kiQ4vHNSFDUWKCqMIAtVsmvpK
4K+trWO48vPYXVkvdalkVSW68BQ/426yAaPJ5sU3kwHHpp9zhK1/jYmL5k85Fc6GPNWizAHgOfu4
/p/3BkpMaoCaPNGwlLCZEbpIBE7N/Nk7bGbbCRd6J+tV7wqM4sjUObuX8o+dBR0LBwSXoS4AvSNo
R6C4UnYKyPg5X6e2BZBqFwx9WfWmxEAhRl2wBPYqDd0kDWtXxxYrH8q9BEpt22RMBWxAR/+I0hn/
Y+Cw6kTxcgTZF/rpP7dwIlNT4btusKxnWMSyl+DoQIsJnGfH38WS+kU8J4thWnJrcZePHh0ETuGg
BbCFvgC2MHd3H9pw84hjNho2ix4cRtUi1nGpy26Fo83e+KQ3RRe+zE2WnZn+m95CO9U/iQJ9fs63
bzLYq7Oo46CjCNRuvutn/RKgqULv5xW13GGxkf4geVsCjTuk5SkjIkUjdhHx2OIa6U3D1M1zdK6H
tsIVpP3TpHI3lveFuXXGx0l4gpT+UN54ZDJkx+gZxqQjROA9/xdKxlsVhB+8Ez6JzirHUt/RgutG
puNVgu+Ut0mlUv7qjCo9YA0FjcDrpZb1W/TOQqH/w6fq9PX2HIcFGlrNbwi2r8dC6hAZLADm/7uB
azYYK4AOVb5YEXmBW19v/o9JAX3kk7h0GMVzLo3OLeuMoZnwntsjvLSiHfAG1VrUDBT/ZIqP6tdP
30/QURX/2WeIfQwK73ua8GlP2Z3G170RTn1bNEAff63XJAag4oIZdo9tyYLoRJHZj1JvU+6boK2s
v0Qb4Bj+ig+cV960xzp0RewVMp2c4tm0CGZMAwKLe9PTAoFqy5+pNSjuHaQX9Xl4u4eBYibQpgIv
S8MgwyRU9m0WC5r9NQvUccJAIGvilAHaUuV4K5X8n0LCM+jlSfW1Kqyx9LPrONuc2wjJia52IHn/
GIFNR95/ajx+fLboPnbetT28Oo4B4PAjmsaoG/gUDIgEEVdX/Ec3QRrDq/Be2cSogG2aRpXylSQz
y8QjwygbLm6BEya6qK6Ze1n/pO1Osmo9bPdja8rkq7WZMluAHKv8hTp8FqduCPDNltBcjBlCeyI9
lgxjxwHOdBUYFKv5lnznX/HCbtShNX1ppg6itIuyt46mXx0Ec+qptMjP0KUmSP/X/MRqp+BzepzB
9VAscfj/T6ed6WHE16G9RnZBeaJ1DeAmUjijH1EEtFMK2kHHnkFGBmY+iZchy4D8DdyO6jbH6ASJ
SlkfYQ/C+RCfJ9Dxla+tkBB3LCkeR/5dPl/9m2QrpP0eBSkhPptPYiJl2fL2Sznz4+nhQ3XoxAey
eWDUY0WwpZ1bmuPIvtPY2+bRu8hyP5GnRlXmAF5xmIVPvQtuSlykfwsggInbJY0ZYN+aLYVSRMU5
mEZXhaNAkLR/SPDLlzC0jfhmvH464poiKrr4LOERb4H5lEHOt+vcGUqzjHrOAj/x34CopF3r2SXo
eu/mBm2YxvVjD3KJaFYcRdEIoWEiWyFtJqzvVFxg/pwFJICO5XyWKmJB2iJzUCX2j2IsQSQFdAMN
tpY36JHNDnfgB3g34XHsQxallKS2eWXERbFSteclEy1YoUqhfTFbHkdV2eZf6g8w5fFHFKUyo40s
30w/nE/5X8XspI02CGbkPiQHrH152fJrxhvcQOoelfl4GzAnjbDQ8lwvF84BOw7fJIom/wCWBV/2
vIppDwKwxMT5vx+6ugPBSv02DEJfFCjRJAxzrgG0k+Gi+E5A6XUdGNMIki/suVEyT7Cz4jyYb7CH
j3mizAPp22yi75wdW9NEX5HvgyuDprt95v3dlOba1u6ZOK9FoFaewcpKlt0lPf2j0tYgkpiWLzVq
vVP9C/vxWWZlzbrXPculCiCPCh+DBfkdm90PaDBCtQcnFllw1u3uvVN4MEJJBHrAv3nWTKJzIHsK
/DMcZfSpbS0J3XBFNf3HacCY4RriKUlb2pitwqubKhklBgfn84cZdhAA3QxzjbvjgOVY3UuaIjY5
S8tMlfD6RliUntNDr7d7JUNiHEO9C95eCBo5DD5i5eNjJuGR5a22H6whAbdQn4MhTVk70o482DNJ
imLo8HZMPDRgpZGMdYy22XkljqKlHWwK4h2tmcoH5xigsjZeeeEHcghoPO0D1ACfSQTHIvZued6j
jcSM4+oUsSTLwWfs94erFJc5hSQe59MLaSdCeeeIrv2Q1QKhvlIjRA1V349XlcRoithdaqCmDecy
9A9+RjVFfqQJA6Tu5riR/PQw8VePjLovm5Qm6IFyFYj5zIOg/7cnsJxgYbscyNk8I4p1EXxFGqjn
D6gYro24orfp+zH0YfMYex5oJeYLfntgUqElJNMXzzcfnDatuDdlVgPFsF3lrfB2gokSpFLinxbW
pQh/hIvl/QsaQCcv9tNFg6PmbOp0NT5/hJcKGL/dvx6TmP7foGmLkCboWYUbU44G3AaABf54OU9n
SDXQS2V313U9bZHVnyaahGoOlzPmvxF9TFhYLRb4HYKUfCgJQ+3lN72pAPQgtTDnDZUBUWH24nws
GW9YIGJGQPWDctMAx84he2v4rLXZf4lT6JXRoxASX3843u/R+F9toNUUu6QZuPER0iE726dG8J+i
ufDPtbxWGZNfv65JnqbUxTaDtnOubUbgBMgoH8+HCoPI86ao1rovkA9YfMYZyMg8iTIQt2xAoBlZ
prc9VIiJR8reaVgsTBN2quQ2jteqCsK9WWeSoHGCMk4NLU7a+HASc8asSSjF30Za6iwraf80ne/y
Rc/60qWdoKf1+dWALtx8MU2ESFJbysXEtgDJ3akEw5UE3z8Cqgc0TrcNKJ9ahzM08zBp8dVRaKLa
fpZskM/kFvn9CFBQsOvhrJ7AD9xeOOollvjI95MsGbDIyFNlbhoo16mmoi7RJ12UDGkiJJNJ3zBF
P7iyemf5F2V7E+IH3D8u36VccjFUVlrl24oFp3G8Mst+k3ZwbIgtSblh66WyE8a6rcbeUMqE9+vA
/D6kH+aO8KTy7Oj2tUIB25sFfElBBW7GOEKiD88YBkPQ7xxBNEatzVkajm6On+JJplBCdgyWC+0F
bFGEMUELob5W6YA3ooE/r0JbcEgjJ2gdfHG+D3KUKVFFS1vLDqyX5CtrtNLHoCWa4xwH6kxiBq1a
ODoV6r3MWBWZ/nvNAhJPhI+2rU/wN3oNybAlsZhs1q5nFjr761K+Bj8E8GRzHYVwTly8Kt1aslwi
V+PNUsVxDNkEHpNkF3/I95lgF4jVuQ+3rISKs/iUXIzC1HxNRTSyLY9h7T1FpeQ6G7CR21AHo50B
88qAAUJ0csjqIr8MQCbzd97Z6sT43T/x38IgsKoGtjiZmyArzjekLqdpJ2FOprP81O34+6eHbIg9
aBj5KFhxw2OW544vQP3yA4mNAlAurPFTGJFAnXMgiXO45VMuzyAp7n8kdfyQC1NFl5bR+d0Y1k0z
ZFYdMJx7tIi589aLqaimknr15/tLn4LbrzgXhH0fWVmDd9fvDHnUBie835guTkINqhVQwDgp8mDe
ZubrlmPUVepcGvco6oGtzalPBCFR7HeDOp2KulazOHZm3EIhP+BzCcrH0rLETStSRBviGhxMOgN8
/m6i2qOuk+uwxH5r50YptbFxyxgajaan47rT5yNdpsWK7+uZEuPjORHoMP5gyMTV2wSFPd6dF5OM
FirdMEmuC6Ek6cETVwzNdEkfQMbUbSyVt5XhzU8ue67wlQA2jYka3Qu3qOjaHZr8LfanX1bgf1T3
W6TqDXyDtqML94bgWSuzU0RoAWoKf2LIlG0JuFnMPaOX4gZ1XDb/A8JHiNCPn2+Fza6rphbUfz+D
Uj4MVK3xX018zqsDT55o2e5KHuS/127T/BBHK2VevX0AA26wHKTqApbdvspY0dVIWEHazl+IXJq5
NjJpRbx9dVLfMBoGBr90YORmneNMSyx25HOLUdEEj1LRJvZzJwCxVLe2XoIlrEGtL0jTOSZfVMMp
3UbdOtnBKNZNFQNmbDcRGqt8sdSq8DTkmrZP+QEtvtlCQp2Wx9YgVXIkOkKjSL2clq8X96+nIt9S
cxy89CzztMSV+eNc8KnjRdhck3+TAy+d6qOz+M2ThEO6CNgOHFGnt+B253e3FTXCTyxY+nCg1pQB
D+vrQpxlQ/GDWUP7nSR+TFbnVOZHydmIbjirPLIVUE0tw9tj1/2cKYzXZqFLgLeHrLWaIepIupVW
ynvEQqCmJ/1hGdvZnRRcQy/0N745siJtUMpR4M+/mIOnYWz9fOKRfN3royjkx4YAOknxvV7snUcY
lVOJVBuafAwLtmczR/pwNIGIm4cgaA9EWBXwMFJ4he0jiqz5Xpaiw6jWKSMhd3qV4szg4mpCLWr/
auif9W73b9/DTevOi9VqbfHXGbYruoxjpt992fhNsJFElx1blkp3fpSf6xa+4whIbqMInOGTX4C7
4ocQAq8ZYhm5x34PoufTusQS7aN4SH2P9oBRyHIO9YDZJOqdD3VQGDx+bnFfgzeQJlMZGhOCPgwL
RSpX7gKmJeNMA6+lEvBCAVjlscQISrzoxT/k5N7qc9cnI/MjTXtW5ZlimFix3orpAMmJThW+a+ow
xdlzuKu1UfDYcpdUfatvDZhcDUa8fVsMNNAhX6JNPJKAO4tYmLzrBv47ltcGAWQLjBpd58C9yGiI
Aeo+4QbIYCCbRiXtvEDkesTxqx43XVFMel5EVb2z2q2+nN/ntwEnCXmSxIQh8QUxTr03bPdURYyX
6pJoiKvc/TZ0G6/gaExMzPih4OLllXWhS/zaifkvREax1UVmG7SB8gymlATmzYCGuE75yW2ZIAo9
ivTY9c51vyMcESUbJDg6xElmNa95xssEnL+OLEmSmVUxIGOyybgbQ/AnqLSl+rhDhGgKiMI49E6G
sBXkMu9tUvCsRAM9aypSVf4w0hefz5bniH87yedzo0b1xqyFr5hXPo4v+SrSZiZQ/KIq4TzFg9md
+NxiCZEllwM7I/yhRkwFocvrwcekruKF0tBaiCA8SrDjWGEusC3KIb7RDbnqXXOoMW4JAo1xT8bR
2Phe3VvDbPba+8+LyzpdcdJNq3LO7RmJfQUCYrMGuOYwr3nrpyGoPJqej+vPs0bBw/gE2AIqtFmv
/8+yzxaTcOIneZynxNHpj0g+Ow0Exal27ol6E8W/IQ40f42hSbCcbg/Vl6OMhJ8Vmmnj7hrfiml/
vEEPXAMpkQ3Uwvi/k5rYpRmn965KyweBhOUVHkDdFMk58bk47rF/ItVpbZgi7+c2KUice2MR+f3S
OGKHbXuZ8d0StcRCezQVgSkJYLAMkvsyZJEzC+IJyj2igP6I5qnya6KEKeAInwI/Xq3afyj+wujb
r90eFhEfjuMbmAlszS+dXuOFRGw0oJO1cROY6W7nLw1CXlclhtuafxp6p+iA2VhjntMlKb1DV8t4
Z6NWHtHPCnA5Z2EoXFkfRibMwZWBB/TP9H+e9qLWDXrwn72kMX0m/r7tgr4rBrAlFMcY2A7OzUPy
6I8HEnx5sYZJg1qiAnvDsty3t065dZ7DFbQt8vw1kubMywSXCOlYnlTfZb3k9JztPCrXWugSjTY3
sSwvI3uuCDJ9tv7EiGsdw0n6Ngr1V1r1+W7FBW5V1sSR0SlIslrZwdzEkhOtlsWQGQ3k44tu6brn
LRCSGlECIrFqoTXx6ojDX9e0AIwYVKOluo/AfgWGmJNXEidOWAJUx+GgFlzgTm3+MK2CwAOvDsff
VLQTrcvdFp62q/B712eywRIqNYn/8HlA26a3ShycVSCqOWvuk1qB/NsP5br3lbvMp5BSLqEZN71i
bMI3zTEqLf1YlGmJXvwst41ykva5+98p3uO19e0V+9DBicc0Zy1nMQ8tgEM9jtadWYZ1k/NnzMQI
fJ9cNEUYhMMpSZUqBXMj1Q9IS7ue8fm9hY+vkWusQy6IbhWpbcqL7ky2ON09Dd3aHg2LBnxCf+Kc
zcckQ4L5iQnwnuKuK5HzsIZGPMbFWh1hjHov0h3IXNrfty18QmbPnm/ATeJ7JNX5sOghNrX9j3IO
rqyYgDZttQOEp9h3YWYTGfnDeidrNYRDcL47ivtFDcuy5zaP2HcESCu/N+3WCcOI39DnP4NPmXQK
FMOjQutk4lCZ+UxUL+FKfuYl5EWIcMO67bECEvGronpK2G3x4KaE0j1hB6udY5/XuCegu8uqAH0N
GmUijboxDhFVshYUfbjUcYXzpF+az+HYStgq3zprzWcj5iNfyFngzq+UPYSwvEaU4tgNB/ucdmoV
Zc75IwzKt4g3KDKzp5iylvl6AKYw9MxSZJ21OJMWtitp0GfQsU/wt7vnfQmwU+8BiMSryFcGErDu
j8rlAKBC+QAi9F+mDKRxi/OF/dxvPFULj8bdqeHiD7rpMrUNj1HuKaWJZjaWmuB7fX9aiOTVP5o/
tHVFSkgXerm1P3p9TMqtIsKLo4j/oi4BUKl0YhaPLv+ArmPCagAwASGHGtFMkx3Bysx5pLOymnq4
5fyaPCJm2KJadFR9SdFefgIa9Wd13fOo4WdecrlPgNQYlPkqj7BGiWihnVGC5BCL6EWh5az7qRPt
ny0FhwB98pYFTDndvH2hNJkTnxE3VKgpdkqyzjufcQRRlMl2PC1fZc3FkY50NilEnSB+9vixCJ9n
UWzbxhA9mLeHJ6V73qJAxF0BrvbDX3GkW9zQbZc6GYmbTt+C4m772WFektq95TTm9kSLbWHc9VZT
axwtsIyfa86I4lAuKnVlx4njcf0E41gaI92UtHA67ISh+Y2Ai0UzQhsBXb9+AIUhl7qc2byESyjN
DwUz/5mtEnV3icyGEtw9LBAVWdB7E1z3NzS+cEt5HSVo+VSf/fag+wWReq7NYwnKz4rsauhiSiXH
ExfjxXAQWS0v1j3hczumXMFrR8eFLCnF2OsgKfFBVYut4nwa3CUK+AUqTLS/Cws48EX//sHMoEiv
Ytav8neciCGa1tey0+5p4+ZpDZRxHdAycFYz9GyNJ4Bu+4jeVV1G3CIb185qJHoi5kaGe/6y6ZgR
eW8BLnXIVi4i7lmD4+w3i+ov+h+f638QQEGLN0cuHkvxiJzcE51TTT+awo9LwqtyZMnuvG634Ius
KvNts6U6DD0IPw2JRaZ52uO+gZz+1BUKjtUQmUS4TMdmqGEjzfQkAriXxQhjcvM94oqFTrXrCzRY
qs797Gaf2Eyz3sAdnVIzPdhz70sMXsSU1X8/GxRdJF35CqNt0dpuj0E8Z29FaqJfW77/KU/LdCOs
sMGQ3tvtOt4CU3w9rAcPjBngujhE1+qjXO5jh3Ueu98yOHCt9vCJPoCuRaWxyYJf6+PUo49nMn4G
mSWmsBocw40jLQp0hHIY//jbi5nAAJr3qLHoKlI13OMuydfiv5Eqd8i1ok1yXGdCkr3AJUHEHRzE
28fLF3+oKayN0G3jeDnMR3Q4ZnJxfVv93w4CWyAW1AnnddhxwvIHKQMdjYgZwDfc2zUi1DNoLeAW
Uhnfc5k9gtxd/StbxjWO8tEQMKlhuN4KnnGDvywcArRRm26XUpLe55Ud408UyL8NHIgIdhiGEfHE
WC7YahyCzZ6yNVCziIG+qyTe4ndaZ3rGOayzC7qFxke4ZNZQUH3GS5FbD2VgENLc7mfbfeZ+ut3t
iXUs28Cg6VQX15DPv24I0kDAaA2d6B6O0H3Dy5/rrPFSDUaWIKlNFV8MwxbRlvWbFkTMYpaRgJa2
phB6kJSErEJuv3BvjBjABuv4lcBcCQYuV0B3MGc+eSx8+VsRB7T59EmjJFVejnqonOUS3Pj9JM/T
Y69FAlYdpAnnlqeCaL5oKjTD4go9BOyxX1fzzhsvsJhswZkXADqqzdflQ0nsPDwzRKepGv2iaKeM
wDq0VKQH0WuSuhulYvQ1FcvXsPucE2pdwFB0fzdx6bOBsbhLI51kD+n/klgxSIlejbo3P2sdmlIh
GIyqtThwr/ezoyazt8R3tWzS6OUrBMuHV0rFv5hCfwys6zAo/0C/1bEIm06x2vkzRcbIGI/mzmSr
Y29T9+ikA24BkH0x+PQeWgbT5EOGGm3cSJtihxDzGEogFeYipNQ2NLBTQS418r38HjzIN2gbyStT
0ZYVHOFcyX4VScsj/5pFM7dx5fs3SjtlhrwGW+olczbeiPXEsMeKj5pc3czZfHT5UsUnAVYETlJQ
DVjjkRlRRYsV2uCH75tc8/2XsjTEjTnuP55L20XyWsfNgKcauJFga5iJ0J7Cbeec3BSO5MO1lbMV
B0NGzIHdvZzsTSz09f5TAeXVRx0uE3nPs/4a4t3ybiewfYZaBKUE6ApggGkGyGRLGgCBtsnQx549
lT3Euzc4/+QzVvGAFciPVO9GoTM2gSknGtiSxoKxU6N9RvHF0pADlGIp4vcIWgftnAiQjw3jQ1vT
XMxa1TnT1RLazInzGyZw0c6Jsrh+ltnV/T60k7plTVZDaiSnOgA17oZCdW6charZHagRVC3a1tWt
WIDyMukyWe68VTaWXC1kwNnYD+ihWBWGoWNYwWgJAw4eYRs6876d9iitFBFlqKRTEyjOl314kAm5
dpxcJmhmTNqtJiqR14nzXX3ig9Y1b2WjrhVQHJYOjlGOjLuVf/nW7hJ8W/YY5uPbo5mDk89UKy5i
wWUrMaZ7L2/pOVHpkAg9Lyz0ZE9Ek6tx6Sc5O5TlCdDnl+CP2+Ww8vpVxriMrUD4Znc+h2VcpUSi
UqqvmUDUCmKW1bdH6WekIvBOYiPLGObf4qncAnRi51fuH2p7GA/aHCzsWGWkevpzVPhGNf014yF9
eWpw4jkNQLJhrKnQk8VVCc52k95yM+lsqBCH0THmYj2JgZhHAClry9RdBm0Cp0BVr6PqwWQKJ6/o
uynbC+JVp7hIbI3NnWMI+DXGGeGPQQCqENcQt6jTKaMS7FggnQy7r3cG9EKfMaqRNAsCS1fQyGRC
SMfPgOpTTnQK3kVu1EC1c4SQeqjBLknM+9qrSV436dhTaM1oSNz3j1BG8B5aNvXq5oi3i0PKSAtE
6lWVDmH4OP784w9XYE1slq/EpMfcFdqEqIXWmgKOeb9SyWO5z/lpJvdVs4fYldNThbshA+35xzN0
kuovcGmGsHPCaTmvGYuVdaCYT5p09DfNdEfTZqXR/wtGS21zNSxmYw/B/kGRQ1rMkoCHKh/2lU5/
5cf+MAP7dYdwQ7NvRynsqB8yzI7l2usZ7jFGVrS+Ye5KPO995LgOE9C/vFdDo45BsMjtY97dAs/U
5Kd0zdkePtPykTtvQLo6G4GkOHln0R3jTCB0QaT4nPvvKUzoW3zyvhTh05On5fkBkz87S8VBWo/7
9PG0pVwxfW7Wfx30iXPK6DiOviLJh7R1nfaPbTx+kEzE+SD+FtyyBJHND53TJT0k+Csv9hNUDE9A
PRcdgISIheynhh5uRgBqmlN9RR1C8+VK1+zCHT+2CSJXrDlbnijWP14Ko6kPwwlRqtOY4OFYJf6p
rva7c3NgAnW8qRyrbnNikKxmubHrk5rVAZYQ9JO6JZ0MR3as1q+PswDBi/S98XC7YsKAEd18Hxh1
JWce541uEwEYamMxNiku36EAV4vJlSaACSCaespuJWJ9w1qWMKjph0kku7kND7hH5oVkJ0lxetCT
PbzY2uFmmHh2HwFbW3KiRKmlWU7UaGeenSqXiYNaIvi21ZNldZspCbOtigUkkHryfgZzbIgW4Wlb
7hEEMh+WeFVW/+zh8rnCDZc526j17PApUfInRM0pdfWarh8f7DYBdVzuG8uEa32oveMfg901XWfi
rmO0FKSj3IgSoY75+xWcc+ZTsonOZvu9ArFInfWqiOXzR/TuDxwvMvw35VEBsAtap041bwgrFLwV
fXg0E+arb0WQSQ97cLSPkdC/cXZcmxE5501qauNDdMNSiHCk4ZS0ucLsgG7yb61FH5OTw1r89yc4
OSx1+Y4o39D5fdabGHhCM6vZayj9+HxRgaPuaXNIusPT4SUQZTzjWmJ8HNJ5aEaKUmbQh4bbhdg8
60FpcFEL3uDSTVITA9VheRUvaVj6K74G20eWw0pBhZysZFmtXc8yGeJPTWxObbiAWXE7JfMgiy+R
RQkjyaKNKtb2blbIMpRr7Tlt6+GDGon2rhh/SNbXdlakE620nKPPdCJaF4bc4lAQZtOKfoowNcwY
zRqhCWr/PRLvgNZk45AGjHOoYPP4SmUIvlv8RYznpOKZmgSh5RbHYcP7ahCItKHSQJqKjHhAImR+
0EMAX0O9FRhY4vze3pt3N7g+OJTOQZ1z0gX3UPGDpfuPCt7sFprMxa/4endVmk3UgDi5JkGQ6A7p
hApp/J3X3BFKx4kwmWvUSLpNnWUUz+jAduZhHqh2r5+W9VW5vXKpNnR4y9WsltpYVZoat7ILmddX
+iN63Jcw/3woPeGd9cZRuH7+TUWhUNF6Jh/STLi1AHX+svS1JCfLYPR5WOaJ24rVUnDSd7cKzug7
w8i7lRDL/FMlb9heAC1x+7OV0u3IF8Meoua9Y9NlpcCqlas2gitQArlt4LhpagDZQFeZO3brAbLk
rM89dbOE9xNiafFn4JH4QTSNAi9lXa//6lyoyuEUJYUXQIqcdIlc+UI2aqyuaRVySCh1Po0s/DhV
3Wjta5z9X13Q8HGQwgOLdZk51aIkDyHNxYHu/JMER0FhHq2Uud8Xo8+i3Y+JH4dSunmxw7p77648
/cAtkzZI87PVWBoYER90iljvTmE6T1DiF/ZsIT5JiUnX02kz/ePk9UYg97FggsmkAwh8TlssiZOo
za5LfN5a/o+PVkXIHkbPKb6Y96GCeXyva4JrXEBeai5ocWe+hwOJupNZk2WhrZwqv/BiTIk0N5ym
ohlAcKHQNCj5G9vbd4VRsyZARncN9H55RdfZcT+K+RqxqKbp0ccF0RIV2R5cMS2TQkfK8Ra9F44p
DQLxacB+C7UnMoviFLah9IW+9lg1Ot3LzV5SPUvQiP8UI7plgO77ZO8N4zIg4Bais3DKx3pEzJk1
xixU5yEKayCXwyAczeAThqPnxJ1Qvkps4jqeCNCQT3o9wS4UCUi66qpb73svSf38u6OFQOxwJQn9
9pIgpToXWezeJr8WAEpCGHiJKkKTFhNg9nXHwvOx2Z053G7izhwTNH9eagqGx6GEqatyyoNanf5s
k0eoOCiJdUOWabkJxGESf/Kzn2wmykaI7OHc5F53XXihpDcxRw8PXulyDFvQDlGf4hePVnvWavVD
0wh6lc9UvGxbQBnChllJqbwTJDU6bu0QzRkHuebOh1NhTKNeBiWkygkz9pRfz6lni+E9DS80Fn2C
sgJvI4lrkDdARgHkmuDtUz7E/o2fMFyBc1m1lREGfAfwdRnT2TYV09Qt++m+0+cNLT4pNOnU8o5l
FHGn1qdnzkD7mSJkzAQkfnQoCnOR+JITJmKCabw76QcaTFrXWoj54AbRnc+xPyxH2kATI1qyG/K0
bwtYSQhAlASpinJBwtSTvnByAfi42xKeiy0xmk+UfUbIA8sToQh4CSmawZnukVOfJ3/ImpfyEBX2
mTGdc3nFK6qzQgLi6MX3aPxWNVLBp/CAfpnL6RJEUlPl2eh40+hfQkj8JlIIj/vXZF1DfXcDfame
j3MQTHvEjRiTkfjcuS4V8ZyKN7U5Tlt3xaUnbdHwgLExEtH1MqKmASO6QgAkblrEAmpY3vnEHdys
asMrB+bLXgk2B4sz9EBxh+P5AgPQ7pzPlEgTXM8Tndi8AfVNlepfa1GeyHtKzl9+BfTZs2VQLDaT
a3YcLvRt2MMacdKz6GCJutBms1ek4ib2SS25CdA+sPAhWNJ5K05awmF20DmME91T/ntz+74sNFTW
p3XohYK4/14p7NVktbgWLJ7/+BgFv95ZsA5Js/qDkypLlyPsBx1rtiLCxkP7XxVlGfWQB2FL3i3D
ZLQWQXTeEcpxA4eb8UonXF1uaAj2oQ77XekF0719753a6g10TylvOSeId6Fj/bdnTwDy7CNb16hw
WFYLy5+ThwPkh01aUXF/TB5lxN7u2SubYXb8lDuL32bujMjFcP/VmfuZNeTnRmAZWa+xIdRs1SIK
QDoOkC/PZi66O33gar9TpMF3sqeSvrerL17PXCHfkHRou53+rz2VJLWLuMrECRqggueAQqgSvNn/
N0yNjWC9VppMwY9zy55mcCRQzIHL0s2XIXRyQ7MV6ds7/TnI4SL90bNh3xOZxtkd6oTgjgdwvXwv
5ZUfVcrPrAKtB4oyI/S3qOZL4Gyv3SCirP07Ezm2eVvkqksQXBu1xYolnqs9oKsg/HIdzyFHLmSS
vth6u0u5bGJEGcxz5nKVqSwJHrileh6no+6v0EVyeGrnR/xh+aMlkfMZlt/+V2OUYT6ZNEMQ2IcF
lpHavd4thLUrQptEVaKDl0+XMaaal7YX98pvO3IC3sheoavWVsJEUgi/F/ytGDjMTQpTCs5CrO2w
QhueKeZZT/cjWXiETS9GFnRo5p15GuTDRLuj+rG3TRSXCmEoexJahS1cTpd8JDrGGrKb8sqJMv1L
Rtf/ZOf1fKzLkOL2DJUvnZt0KxymJDsl1RX9Bl3HWSTvqyb7pFlYoc248rkm8u8LsY/X91p5H1oY
oWbOZ8fFuxvvlWJbJk2vWihz9SkPvWLKjzI4a+vRHLgdUK+Es/XJlx1Not3QykTgJMQ+madVX/wX
Fzxxs9/j4fzMT4rES1Exl0yqUM5ArsOqx7TDGK/hfDfI9+8Ttxxu0tNkIYL2V8tAhb/r0mR63f6e
2w+jGXLVvTYwmU5T9jT3gbJ79jkt7ZbYOOBqS/xGlvEOM086EJVWF0L12Ihjq0RaWq3UOWyUSN1x
oxZv1uFLvRJZLl+o6HgK6AyfgLtJUJsse91aGW94+w5W6pZB0bif7Qn8VXiNIrhMypncJR1sq038
iftH3LB8USiCmwpBEiLkfOBDHTpFjIMbb9HNf8ww+5Qa4fHC8YPdvCsg4qW2MqvI0aetTvWgd5fV
TyQ7nqqYGj1unc/VxCve9HORSYsaXePJ4rPdPZ0PrFSXOA+LZwo0lINW+sUfQ1mdZVHYHWlDnWEC
RZO4n16Wpe42gQKHHdAWoMeJCb9kwlzU8oCZG5jvsHqJZ31ZvShNKKqVbLY9oQfdqkXsj1SkIrcf
SZhfEtyGiMO2s60xPkUaFo8cffEIksSDFJ6MsXNmUW3M7h3Ejzz6cz5ZoRQRX8ei8g69h/Kbwb8m
uIkB6vURgrZlkBHN5zcE5C4IJ9KBV8/wUZyLH+ireRzlBR+5rZK4Becb6AJYOj1sAPCSnd7i75oL
KvqUx/nljaFscRu0ugnHQQb99bJBw6TYHX/zy5T1ur6WGDnIbSvxV5+AuxlOBYWk6HRrolFftMc4
jhZm74ewea/oAisOQkup9cLWfIZAY3SHAqh+uL3aIeXHJIcm5yvDRNpQoXzRmnhZFpJ0KlzadhGN
dxxrEPMZkEtWE4Wl0pqbBFdVuvpLEU3JzwqUC8ydSQUuv/0qVOMdJ1hU+NFyRXBU72kK5OLM+n1M
KM0PqcogPs+/l529GaNSgZX9FMK8ZDWlAObfVoKbxayPkAIDLtHM5nCKRrHdoYeArcbVY7H6JLS+
E4ge0b7HeRT482xurPobHIQ6P4yJw8UML5CGDU5yeQfwRMUbZgPzbREykKqwXuG+KCsYPckPAgJC
FmtH2mSz98pu29uKAoxt03juIac2RzTOTv2tDCJY3Sm0K6P1CQ8ab52YVDAiZAxxF/R6OCxZdCR8
gwXlCr6fxq0rYMKCKyKVW2flxqbmVjW7v7S7ZUVWEW6iIVgBnEVmSQUlUc+0tIuC5MPk1pb2cufL
usKLd8P+VkfPvLM64hrC0gGEa3KEY8bcxbXqN4pkUDS13BNHYJY935yKAoStThchP9EwVS3YyGRR
/7UiLh87HhofCW7px5swnB8UZSOUn7ZEVkmi0l0Kq1Bx62gtypO2Mt7ixh7LPBkvDE+tLnVDmL4J
ExeExrsf+0ch/NXjEeFeUWhJVNplocHT4Q3lxos+FzRSas1ShnvpNegNuI2jQ7i6Vhh+ko6o9Ld8
swnRoxc6FR35ch5N+Y59JfWaGBPl0SsuFuGdI59NWSmksV6wDsuSB3jlJQSLfonwnFI4Ou1DCc/y
rHSGMM34SvIwAomh6v2YxaE07Ngp7RI69oifTXhPQqHP+9VD7TxQbaEp61Tah5psWddfzTe2NiRR
3b0DWEngnIFzbT1mGF+izHWEVFl+hm8lTpjbWC5HnnKo6ngBnhCDy6LB8Jonq56ReAiRgXa0AubL
tE0rAXPYCmj3Oa3I2sq0Y5+VzIgV4//nIaaZn7KBIx5mtRwCFZDnXxE8SHjGDcx5Pw1ka5F4wYHS
jvBZkqXbPF2tpshNjS1UW7P+Sh62QXbq4sJ4SEmjSRnmON9W9cnuX1PxYowE6pv089lgqqLvU7fB
0nJEtOTMeEqVdkPI9jX5W0IkKZcIlEd6Dyol72mKwFSNWDzyOLwhzsUlKLf6ieB7A51iY0jpauC5
TerRHPBSexQxm8cjq6NYOjvuA4LHu2cPUgOEi5iPgFMdL+HqMY0HQ8hTXX7h+JQ31btEqcHXc0AB
u70g9P6wpiDt028T55gJObP87a+l7LNnzmRAV/LcV7ifaEBjgrceDXS+/rq1iZvN6K9VG28VxPDf
+KR60Asezqmk5aS35t321Bnd5P1QwxnJCi3hymJzVOkRYQN2Vrmfy0j4QY/+09U3bVqRD3wrCNU+
s19W7wb66CbdZy3JM9WUtwmJQoQ4jWrLff24bFkA15uhy6je3qKlLrEICAQUav0D9SA+iAty/gCY
75SnkzRx/Xfo8ULpTIrXQmVQi6aUuHRcFHsIV2QHVXiesvnWzAYmHm13hwRoHTV1+KBzslkP5zZu
fU/ls3cZROhtos8dNBsT/Jbb2mC6Ogh8wlffMvYNaNzgx4iIu9BrTNV9CiWH4nNnjLN4WD5hxQqt
j8TldwlLi87r9G2K72svY2dv7Ulpcat+7zZIm83CEVIUUoClkMb0/IkhLbP2YOmrFYljyYnEle1e
ccD+/Kxafp4lmqito31dLvMBFanLTpaD/4329xnQ/CGj/HFQyl9X0EVtaq+8vptpILWt2BOex1TU
KXIiPf/tGFv0dZc14eP2V7lgZ9Elf6Pa0Vn8AQjwNsbbgs7Tb3oFNQrsruMbQ9lqCQ7UuebpCG+b
24/BjLAhCk8XGErLw/JGsmPR/wazUhjYHqbn+69KvmEK1NXEEigkZ4SgmrWpseoGHC+2Bg8aFRiO
Wzg12hZkYK0R7G1tUrQMyl5YTwx0BDTSrGanEoY6EvId/JAoiE5bgS5CNZyWpqVV/o/QvqxSZ/Pk
J32bMZh59sAkExkt2NvFnbBOxnDwgANHP0rB2Va8MKUBIJiSZlG9ikf3NYg2VQVO/UGa8GHEBRCL
CiBGFbb0VBUR6c0o/FJXTbeXEulXQlN+i9EJjDlH8DRin9qUrRzt4uV3K0YwZRNpWbvdx2YZxo2j
7v2CqvvVqttu/0NSkIsEIIwSi+wMZ/pERYoqKf3/OJIsgfQt+gi8EQvQOOGqEMLMmIUGyOPgLOXH
23XjcnTQUJd5HMmiHwByJJi1lRPKB7kIFDogLhsJ/sZ3CaDiTA6ORziBa4cjrAVOxktSedfvSFkQ
Y6KSNm7/1ieMP5H0C0qInE9C9nXQn9Jy9orMsMrJgeibaKIH3Z9i/DSPhntEopfaG0fj4FelQVwA
2UheOO0EFjkrQnS3bxhETjmajSSmXhWKbVGYW1Txj1sUmz2vU94tjczQSVt+CSG8fZ1Yv38YbENx
iUC6eLMaQ294MIfSPGiDE4rUoULJ5jEMl51AbtV9fFePRr15rm825z9Hbn6sO0dBDuiIPz4WgyMp
/YtDlN3p94BV3kb0wmeUwDEAk5b2hEtoF5FJu29bQXHZSYbHYQK4rMs4bS22JyVoi2ghSFREE2Zb
Pf2qm9JlOWtsXpyNEBwN2XA0Kok4f6lvL/mNpRX278gIL2wC9yqs4LlF/yox+cBZ3rg8K8Q3so+F
dDyPRQbTvmB/iYllObNrR/ZEl7h2MmY+VbEk0c0C2XxbTp3bfu+zcnGk9rUnPA85tcHKM9ktLO+u
A6s2V5l3sXFUspvu1vtOLbBTLhenb1A888fZUyA7hPvohHg1FmZf9iDM/5VyzpSxW7/aBUOl5JU0
EYRLf0pBYvJxvc6xC7QaaPewef/EYai+d6CPO97kTdGMCePIW46Tz9kD09iyAxV1C46QpkbHA9Td
BRbI8/QPm8/h/CjL74lRkQCcWMD9JIcgZhPvnG2YvFomsTXzKMAy133gJrulf4XxxQlJhKh3+rZZ
t3TItc7X0k+mQulAkjunn7z/9yRnRaqZsqY0PRs6R0TtxOEWW3ESWPWvOdPjEaFAAPFVVoqXYw7U
ZhETYm5n3kz3wSayjqqsftWa9wTC1hs5e2ThQXb4Lv/pG7r6cLZpbf/KXtph1RjADjAokmgPyuFS
XB4wNYWH5fM2XPKa51Ucwc8jlJnu73QMER3VAPHkZGtLc1XTW9vcxedAmmN2pELc/VhKhaeUJlu1
7n4mCHv9yIaUmE+IjZVlQOSRHOQTTkP1kvi5gwTqGRCvDmjalvr9IIcTPiJjQGmVDUrjkfgygdBT
shnOd+bvQlhEe/emAby5bZTyUZ7VXtUaSJV5sSV/zl7K/8xM2GazMSpnRV6oSOJmuLq+m7LXk4cw
cPG4/qMsotBs3r9rhHz1fdwZc0nWMtHnaft/37bk3Mr89SbnM49aAsvvJt6epHWeqP4F3qkrMgkb
lUNs7rEVrJOATr0534pFyMHhV5bPTMO7DgvQ/PPOxLNilAq+Y/+s0rIrEuLM9Zjzbr5WwO9Jhdur
C0q7XlI2JiVSUPyQFRG23XCgrRZA4VGm0ZbKGocaay4sIacCI7tHkVlNNsVsbD0EUaOnhxXbNNM0
GkOWp+3h4qjPNYaLtUaEIv/xh7LiLrqVeoQHNRaS2cZaSH3Se/U2p8EH6hWGTSrW7Q+uRX656PF9
9t3oxJRGvnf+eFUEQkQEQxg2VdT0UtRA2veanOboe7xGCGhjd0cN5QOJwReS2dEDpuLLMWu+P3Uo
eQCkBjCHC4rnJu3goL9qQ3gDB7HLCiJA7izna4NRR1jQNmCUswbScgs1vHbyWkRberSNWN4RF487
5qv+d9lT7Ix+vMY6bBmHZ+UF4z8PGGYSbxNZVcGL/CXGArdeg7GnuCnrAR2jrNwr33YeDcYEmJae
421YuaBp3tJxDF4y+wFliGwk0aLQ81rWdDefEh9nGkKcJl5Zrwo+kRKl0DwJJYRP+e3R9udP4hZO
JTM30rhRQAUmWiAwoWB9VE0H4C/pHJCQRQpAGfFWZXSWWymcOZCzZgLcbuffhS8GuB+3zgPFDhnx
oSN0b4sp0YH/7aRQk5HafRk3FyYWwh0paacSbRaT8gwoiuNFmk395R5HWPVvm8iuzsffSNnyls+N
4glDtgYHt2XpNYoLZZd5/Ej+bwnxRBHGj7dbxvTOnh3IoHoVWJHpriza6Zao76OPJTByavGHrKyO
U+EnrcYXyO9MIyIWewlRtBgnRwqSAA7g7rXgcqRYSL+SfQHZbmHMtaoe1enVZNH/WIM2sUA1e3t5
eCIRnB1N+eZrLVFiaCBAXXU4aq72W1yMM4iUTeD+PYgTfDtYH1RJFRjsfq5CDMeSEHy6gc7F6etf
wReLDVAkk49Oam6gNVtboIMnWzDr9G7uZNH7d3+6f64Oe1CSGAvxxbAcH7nB/HSqh+xnwcUrxPwt
H9eUd08fbB9OfgwxjutGHnIRYKpBjiu13QAwXfExRWvdwZrsX1c3v8pGgVRoQip3vMQ1UTNQAj/X
hGOMdOBKE6SYADIpDcXYD0mf0a/KD8QYurKMRgx7kd9IfKDaCJhWMliOhanPO89D5V5eK4VsgUM4
/qPv3a1gN22CAsxcp5F/lXDYK0RZBJql51j7gG8GQXfPFOSdOL39pCPv4PSmiP3oucojkoppCBWp
0StSWd9qouGmAFPjYE6KzEwe/H5EXqOSOBLohJ5xOmOrAOFHQsjgWkkiNJSTpz4jC1LdDQ3i2BUH
Yf6J/G0+ZR/kcTsjLcuF410yDrupI0/j/Cik3RD1Yqf17wrukZHY/0Hxf+kd10BrH7QcOZM7t1U9
u2K1Oi3nc4UMPm5jkoaSaKoVIoQbgdq6NcX0zuWgp59HyzZdI4tevAHlH4IyFjpcAJnnDNePuvDq
vUkBz+tY3c42JNAuHAVlZDOgcKK4HhO1xcIjm6+1LzuHq47sWqlBefdHfOHMHV4WqrfypP5XcaW+
IyrdSUVoP46rzatsbYTGai5BihJzXSByjwWRDPfZ6RCUf33ByM/GErHwYK3e3HxvV7K7l7wOoIdY
/QkCHbJN9N+y7E2ZWymrua9spbxE0e9glFj9yw2BVbYGJxsV5cjebmwXOLkaX8kdcBVFQovpr13c
es1uivMpoOjoqEiVjcHi7LEhV+dP28l6vKehO8oA6lBHWsIYq54clc4xa/vhSUu2sOedliBJ7sDb
DU8f2pBJweWGRAo8YBndcekxPiBo3PRyP0qVKGcLFCqoyUTRQ88Dijy+TFE0iEuji1xi1oU4xG2t
ItC3Q8zrde0WoaY/D0CF9kKxxcrwQBE1qnMGvLikbBKeDYnV2voxyJV9bTGNQ0s1S4rEoKOOQZat
Ay2iY68qA3TVMLcHvEOLQbpDDE4h17+pZrFBlokqRH1jIuZJUrs4Gx0mpcmSbZhiPfzjbuRT2BkA
ebJxrllSpGJO13hEbPxUpVwXDJ7w16CTQe4sXAA8QhlZUVbuL0DbKtDm++tJMZODhrQXRzJX8cvJ
iRJ270WhhGLVNuIGK7oRUgfuw7t53wy1K01ZcKqZGsecejUHWEQbdfiQXry/DhQa/M5+umFGsw0L
AYx+rp4z/8Cd9kDjB/kwYB+gfUGnJNHggOI8PBAg5wqE9ySLgXVI0zIhWR2zYxZ1sRlmUV/dEOaa
jdh+uKGiE1d/GWPAHqHsdsXlMrrXBvkHsPkQLax9wq9jPIYmDo2VkRiazr43porsWgweu4SbVn1L
cgNfyIvroU09RcLI+OX+vDXzTUTm7T5+D1OhpjTmn5zNMDehVLhmLYtdeqzfmkcJ95DRoAFP7WuR
LmiV7vD34ox56ZnXuXbGL/WxwQejfrkINXiDjpUnMLNSAkHfj76b1NuUZJTfbFe9udCV+cl6f9lz
OYGYiXKWXUE3HTtCt7yG6ussflreWFqaL60Rjt6PSrGQZuSqJ0VrYtPvxNIXL+Y0VdQgrxU4OPH7
MSSSG+knxwPNRIUtpAlT042KtlPe1rwDPi2nz8t6RH9uESl1lMXMGwNykPfd4Gz5TUr7D2Kg92s6
6t18pTJ5qBlhvQR3h/f/VhuwSnCzFTZ5p1A8Xg1gDcF+VVZ63pWJ5zR5WOvJt/wcBb2zQNT95tWk
3ZJdh0MSBJwH3WOMwF1U/B7qEhDTPuLseW9R77h7f0LeD7TNoENLwWog3GBWZagiE6jW3bEq6WEL
g7n9edM/L30Y9wT0oi94kvthVVjugtIwjb0HF7esMKgFXjHQ1pJ6G3UMsdjNsvn9f/CE3zW8o1ix
p4V8xfufzsIhiDqtudTiVXtlaP17AECXt9WVdNx/l3laHLB7BZb6JNvbnntQ3twmhKETt9aboqY6
K/kb2o1oTEL9HwG8TU2XlkiX6ebzRmqSQf/g2YfpP4N2SuvyfoHcp/J2IRI4HZC0GjxJfEHd2rrq
E3z5DFzhxut+IorZe/4yEeWPkGXtEQ02bval9Zn2icijkXKzjorlTWGzW/nqoDO4UcyTJFraliFK
t1F85BmssuKdwUFNjxA3Ptaq/81sUbWw1bPtfQsIILFp2lvZ4ZIpCYTuBQQw3aabG+CyDu2ixfEk
tuHmXiJaj6IHVDQH12R7BChf6x38Rn1RFZJ1Lwb0KvWKVQX/Fu3owN+uv7KEA5Zzeq1cvZ9v0IEF
W9sAlcziEEWDFKox4YDM4TnJPU69cvQhY3ejSPQwCpzZtORlJOoc3faCMMBmPpYNN2owV2XVgllW
lq4fudRfFexUD+HOTwS50ELu2I/kChS333Yf6lpfF4o9VRoTAMamqkOSGRYBR4dzURlwLLTD2PDC
fKzkga+be/mOOCQKEwqAvPnEdKaEQhZiJw0ufXZyPJQRlIId+FAcb2Aaof3ofXrKqUeZAWpF3T3W
DJcze/bDKfUK9I/2eBsOTwzbD6N8G4H9x06fFNdWZr1aCnnFVG92UlOGHRtncbwG0N8KBY2HKrgF
ATkJq0xeuqOc+FVUgMPCx/ixYJxxs8odnUmTecYJcyxLYGE4ZhuP75+EaN0ZfnWamE1zaKpcs4tR
7u0cGi18Tm2mebd+AWXBuGJSlysGZbkVR8JB6POXTeomy8m3jX8CfxT5mgfkeE0Tvf5ykuUVOfjl
6EZjC6E2bKRD/Hw+QA5aZ7jsD/Mf5hskWci306Y79atijJ28JkMwHTGSawatEBl4YJ+jsXl15fdv
jK1YN1TvU+Mto+O5BTfwHp6IjWzmjHm/0x4rar85JVMGUDVR0qr26rBBdRUiwbiLWY5KEokljuF4
MN8qH6ldEhY2XCxjSi+B7VGSC8JvTpc9orv4DyumHIr3lxWYdUHCu4igZtLP/vsWaQ0RFKbRkgTU
JeGlkGwTE0BhUbKkn19Cgg33/Qqefk+e33PtTDLxFtpWmEM8dS8S8rq/bDRhkE4V7OnO5oGKPjXx
a+bF92058857PQV16yjpO9wdVHHfkXeiQNo4tup+ZB+1eERUZm1v4UIILkVel1zbwy43wU2vStcY
2fQgiuGAR2XTzgziqcv/K0gvGAlrhEtdu0SvRpu8GWIQ7s9ptzzjCElNKK5MdJdHrhp8qEZoWyfM
FpzyuvGzdGeEWij9917Gm0H8ZXtZqeyRx3M7q9QE958EYVN5RmZPohwatp4IBR+Sah0OYqW/JNlx
RHG0LRhDVEGQOEXHobtlmmJObNMR6s0ghPgaFOyD4O5Qxl+fH0jEWqccb1chaWAPbn9ay7KxWNS2
HSIbGI3t4eBNFJWt0UYqAdQcvtS5QcvnHoU9S6rv4jKMBSRx3oBAw7srhUpb8EPbBRsJHdreVD53
J1jCDOfC05LfC4xwF205VkXCAJ8IwB0Z/MSofldfxMI7IMkRLPFYt+7TIC3NoacmlbgNDnDWnaH/
nzynt/fECLfYNB1ZPaifVgae9NJnY/h5PMQCtp+pQoqSFI2a2xdxqZJY/MyBXD20lmp/dFnefXGW
DJhbsWRFXpJEWRkaiCsHsAxQnC7ztumsMquiV8uepdbIeptFEGhPS1fRPSdTFpYNZQVbMC5LlWMW
P9QoN4nIGr5Fc9IBW64aQBqGX4R7dOsdGArLb/gHGlTm2ojjr9Fx3DqxIqqjAaUU7BYmVBz5Ey4N
V0n+1VbOTyYoOEC/pnP02dMoWkkVm78BRmurK/Xkc4kH2kAeVVUcBidY8dRRy+qEObn5jx/R+qcG
4PhC9/ODGQYo2XKEWf4w+arUh9MSfVo2+xJ4L39jy8NwkyM68nzoU3n3Umdj++Uxj+408zQc2xYc
zXZrNWJS/jLIZJQOaRe+zAImI3CBO8oQy61zBc8jQRIIcdblKaZe5ISEwXUTDWAi27rfE2KsAbM1
zXlIjaK1mLnNaMJIVvforb8KFATu/rochGgdpOg/EovgLZxazRgTqA65dNgysMm9plcq+e7dUKaQ
fL53aDRCAGv4akbBsJqgqm4enWNRMHSjKr+n+fzgOE6Rzh3f/H+hMn4YJdjZ3RNYuQllv/1tX1zh
3KcWDex5Zfp4bRKoUOxA0/oCr7JbQBYz7dQO20ywBe3EVzOJLBLUlp7EEthyvfbUdFtSgUlPE1s9
sMyWpBVmqlM4pqPhm5CdwywJHTlgHVNOteJGd07m8G5S3yAVu/L6KmkbdLEkpaQb0JrbimvCL+jd
9LmUpwYWl8Evb28zPc0wYREQAv4v+4H7nT7748uxYNYmNtuSVvYEJ5SP+xAj4lpHYzUY04ljEDiI
9PdFD3uYnpprNnB82cMemy93+wRUy3Dyh1/Fhe9iVRWxCnv11AglRbX9Z96O25w7BFw5K9FZQry+
21XRONUM8ZEBlrbR2M3Z/L+vfexMeuZSlPTMxvhsgbwyoMUgkK2T64+3gUL92XfBxjCma/hegpLQ
SNKUnuscrtj7woJaz0GZWE0m/qCwVTEyS/LLcxyCIO3owVepeBo0VtBPc1hXdpT09MAuc2GLkWoG
w1uWSFJhZKSJjNujAM78eLjBo8Q/8I1yjKmnaxBRUgUN1gGkpKNHrVSl2B3GLJCjpdW0s4+kwdUE
085wTtc7FlwHLecyRNMTw4AwPbxZOsUbde+R81XRP+d3+wx4BntRBK+AvpL/T1s5xhUMpUFzDCgC
8G0/vhFCBKymivfOG5pTH4574IskoQ5FU4oWWuqOtPXJDgHAvrBeefMw96SHwjagxjy+OFjQx9TI
gO5LKxHFQTrfHQxwhfKdBKeaZAHbRp9f2LhyWORvpduZKwmGjad7sCbW/9UVQ/6V6jsfGULv+B/c
tDQRBAjHyuYql3ZxRGRqYE/eKxS5vn7N13iVDSD4sHFKjI6Vb1ZkFjPMUnc0mkCxA417cISaBQ9Z
mGc1BDYC0TgNLYd8L6yDyi1lfcuR4cqdLDhxgyhir9u4as8HavOn+AHkLLA/iRLmDLsdZh5e9N0i
ol8FdKFm1TF2w+xx/UZT0iPkwdVOGuyVanyTkh4mJ8PjanK/l8OXLOCmHFXdhFjYNVHOP4D78LGI
68YH54VQscGJEbvBL4+o9vf27jHZY22snQQ6ViWLCj7Oit/KXVmzNnuFjMnIf6mX2zfUmbMdrWvl
2Cjp0hToFx6TzCZuTflxih7av9eSU/NcNMKflxTeOWVoJqjo49mcou3CcHdZ7eWbNg61nHcb/FKK
wUFnfjLwOt1B3u7Zncu3sN1ks1luF+oXaegMlr425885OgCayx8CIuOwDTjGAJH2MuvRC86ZZWuI
5fCKHaq9g9xz8SjHtERQVhAEiaW/DGbejxvsZFps6cEfid3WxVKYI4oeJPZvTIX7ybKuqRdk8EL3
A1HvkVjc73fK9JTjN4RYXw8fAet/Zd4VXFcAD9N04K44npqCFTKgB9rIyQHNMfM9fyOFNg2iAbVl
Hkl03do+7PEssXbaX6240mAIjXIayUCVZjr2mGfn9BYnw6FMWFo4xaVdIELnsGLvD3wwKlGe2mtb
qFc7njIaS02iCQwPi0PJUCIor97EElZ6C0gTKdwqp8kf2sCdNRHOVeSWghpJgJSr5z3dK14kIqCC
XwsxTa2xCcWZVFe0iEg6Mp6kuqWRN+DdtVgNSoZM8fM5hGd0RWTqyuxnz8+KHSnI7de6KxCcE0SB
U1yxJamoZsI8oKIo3zqG2jr3BKHXqUMsU56qOc34D6pPHAMpGUHtBaq8jxuzLAkjSbqh4qwTvs8u
4ccywTquX+oKHwJe7oR8P+Imsy6avGr4+5vwbrXJn1Lzhx/GxPoEJFhNMttQpG/LBfqAfMoTzaC+
Cm+xW9OcfUeHfPQfKZd7P1wOOdHIuH7pnnE86zRglAFGOculs69WM5EbPXAt8UvCf90PTxbN4h1K
lCBvt0WC/pgSVY5FCHAZvNWbbABxp4k28T8Fs+Gr2MbwnWYYfLAxU9lD+K46A4ttOUfO1I8BT/jN
1YAjI6MQOje3kfY+xEF6z4JgJMshylGQKdKurl+qx73vuwKlUy9ZFmXdH5ghig2K4rkW3tRnFzi1
O6ZRifiZ4Ss0IX6Y3cYn1zC+lNawTkt5tqQBRrS6G2gjgAohb+LKwAcsd+n1oQckfZjZ6CFLKfpr
PajejHc1l8BE58CK95lgTxJFIZAMqlL/178ScXfwU+8XdNupBzNKZoXwKWTKICV9izmTky+eBY64
ZJZR/wRONcbFB+SUg2r2kbLopzmpwND8rMAamScyQG4sXPTG7jWfbdBKE7mjE2OTX2TcQha7ujD8
LGDv5bT1EeFiTyfd4A7CVPZ7TQm7UyMrnUlGWYVW0IGfnd9BLafphj7DMV10n+2nlSY/YmyyvqOd
lrWE/pwaS5Ola4qkvar1tvi41jsMJDeYQPAl/Zozj6PKku7odv4NSpc6A5dB1A3iKv4eILGWIEk7
++S1x8WLPiU9fBBFg+uq5dzCkuFpZfa4ixd5m1pa34ganzZgIYTmykGArhyWUFirb3hsnz6zij1+
8iMrtmQr9t5u5tUtd0NUmhc+rzZWhrg5EjAbwFzk/P8PvBG/TmisNHG9+gvzcDvORYdtcpdBnxuC
ZiP/uRNEr3YcAPfGB4jinRXRtgFSzG+Qjp56uyrojweCatz7BNNgB5gszfBN+b3VXsgUEAg2TU8K
yPab8GOuaySrauG4QqJCcZ7LOBd0cj1Fn5pMsH1iC8z9f6Ve0R5/5X143r/mv4FCAiWdb9zRsGCE
eEO5NLSYupbBR/9uLM9S/h+jcqoEsT5LseKmaCK7WjimbPgjfxnOlCE4L+8lKbEJb4lMVinJvSWL
t3h+BwNYzkLJEXpXp6KekVadZQXyOsY6MWtZ+HJGUWTlnoHBQxwfs6DNZQzvTbaC2A7EThFhbZ0E
8qpUpgEc5siTZa3XVrHwzpFornsRRxiEn2fSZR3NfrdgP54xkIwPb+i3eqSatmdrT8+OT1KgKCuX
fGf+IsQnc3gjTjtaYCbBGVKQ7EdOO8sOWCwh32S51SaDrOP78hYhCXAJQgyFxfPjj3QovBAejIJJ
q3vCuQwR9Hp9vvRq7KmKhXxrTw84djHNZ9LUcG3YPHBLbI3RtRPL5sOvxjhSSrnev/PgYl6a+Zmk
gw+M0JJbCVvpQjbPiuQvY5shfv4iMI3PpoeDDlvW8ta8v5KgvWld5ZQr/0dGfB4Q5xXNtOvWTIG/
pLtN2nqCyHiQm9N42X4S6Dja1abVrwkDy23gmGTquNH0ZdpPW3JbaeH7JYEzk2mLMgvgFAqVxcKG
7ZucFv5o01kMGnufhyA5my/IPDkBkBbUER5jjUVquvYb7Yk1csnqJwxqE1OKhzh3BAKlxJL9ijYd
R3z0c7dgQoVU9AmQJRrJqn6Lyh5JqiXd0YUf7PGOjuTf4X1B5d2JReB6qjpYyCIUgsflgE2T9g7y
7QFArl7hxAb8ya9FprfDMqCyo7iaA28lhaRDSVywiZ1tuw/ciamlb6K5qPE6vdcxfE/Bkk7v9vzp
xjwAAK8DwMxzNgoCA6F/vDaHpiSeMYcmp6rdkVPuhXx9Og0UKZ/JVY6sJEbZhCjtrj8WseJX9/Rs
CHUyfnG7PdJayPdVbL4kipgKczmWOBmmXELFhfxtF3DkpMvlBKRZlL7RhdiJk2SN6LIStkvxrROY
3sUhK4kd2ePCY5RTWbTDUAcXZxn7eRU9gT3/tRpoe3goSKGY+ZGrMfonjcY8ukVVKWb1WWB0FOte
TjDo/BXGAlHzPtyNbRr5lz2Bb++hhR2qFR6n0pZTlMkKE5HoU9TX+T5OMG1oC+3J60q5Y+viwibS
wrGlcyYH/DcZTV4lgq3n4hZNxeMzcVxiUGjWwgCkErXp3oU7OI+F5qyKlQ4IaoBkQe29KlLkHMGz
Pwr6t3X81vrNNEM9KqXFOzzyS1l3xtnFht3Fwd5OjufkwQ8nOzAWm/BcjR1gFeMmqa9EIiRycLwf
popuvlftM0GhUGi9uQ/ig3bl0RZ2TxeUaS3nYmHWq6l2f4xqWM3xWe8WpzmMC6Vg0czC9VKIw1nj
Ge4jaBEcg3imnd+0pT3kpgl79ybQo37RwyhGesXMIrTskmt/qavBTnQTXzUtiFRr4Ey3scijJAlv
jxGheKuM9sw3Bkfy3Rq/k61VlKaU4r+nHl9i7t4vWT3yiIpLg0/HOSSumLZmw8KeVDzeiDq0iWYs
yGG5ak0IhdJHEP8kxRYajpqj9OajPh8qUUJISDLBU6OBt3hffbl7Um+7AVRlEHJH6hQO1LYYQgXD
XKm5pjYkQZYZtYrP4Hdpf7STtIHl1lwJAMKgl9J+h6YqX+aLNKZm0YvwZ5/iBCJlfUqD8kACKn61
gh4/+p3s1sxcplYKVT4mNWxUs1fFftMUWTA7gfwmffMbPdhURf10g/3xTfusnQbl11axM+7q5Abb
o3s6jorhmAHh9h7xHKYErY1kt9zu01B+/NhuGB+qSUFkq8IhzmjdYURvZPZxAN/+YQBgQPPV71nL
POpxuvKq2rzS2pSl5XoFY8GqyvKl24n3mYeZJKe4AdT2zbfF1pFUPCMGh01e5Ey7XIQV20LlMMcI
4oZXxBHcqqZRqu0fPrrHR5oAcPUz1ufms8iWETVCYPBaiuK9aoF5h+hcHYSbj9kCX29eZwievDeD
pJURRRNLW34y00lgRY9x2mX9udugt9PlXlaOPzuzXxhgFnCxAqg84U3Lc8N031Gm8ZpDqzQIb69G
LSsguE922RppuiNHIJRjVTvx4X8As0JkHLePSNRuGgSZ1ucHuAXBs6rAwrSdd/bsq2/Zn1epTnUl
eC9MT9+oaJ/QN04em60FdAWFneKSc+a2rzj+kGzYJ2fpW9jiZpcFvIp36SwMaY3gYakFoymBOXwf
3dvuuALjRFbOXi2MxthrmwCH7BTZwd+ZtGzHWwGANMN5+MWrn2x/r/6k/WTbzn88dS9Zm6aJ2p4P
vGxWNyiriGPAWY4MLLOVNkanflBIG9aSRry4iVKyv1Sgjk4qBy/U8JflJqDuRGnech68AozsGkvu
cFY2GfrofZLcw1Y75P9deqFXW3bmYKQpP8lL2Zdh5xf8/ryHZthtS/rAL0mYQTW36k9AG7Ua6X4d
oSwjGh7F6KX1bc6m8JA3Td5BLJTBT7Ins8YajDcOgGpbInGRmapLr9raFEwQo/ZPSMphT4u7uSJ0
HnqREAleHZ7xO9Dwb32cfOGQEVC98H/WwB43kTXE/aQOtBn8Pt0QHIVZzxBES0EF4qMxyRzxcvXb
YavskbfQtNRSoJxJJIoKvttC3LOFD+tjtsxW+DNNtJXCmbU5Bq70v0ESu3UboCjZd52nlak6zjbI
+wBWK3izkO8I1SkVkPzf461Nbs9NMxg7A7LsrEtOhuMz1Mq8sF53BUnNU7QlEzBdFeZKLlfNnR8M
lVlGln9NtzJYKz55RSnKWxv8WmVbwqsIpUgXLKOZ25sdvfR+e2Q57oSUoYk2GzPe0MJrXzazyc3Q
D6BYEv82Fl7kSIbN4T9PPz9tmAViThnGQEaYF/lLVz2hRO7Zdazgk2gxHEj+DzDYe7726U4jEjTi
cA8w/NTbrobHSPU5js7avNMfc8x3gdT+kXfpPARO8/FCM0slIVP2HLLbDyIjbZI+sRKoIEsNt+qd
0/HPh0/gwvfUekaHrl7QH24nM0JaTe951OcbdgKZO9xRM+x8G1wzBecH+YzuFgiJ0KZcj3IyqDRc
wuiijrpWRrDWLwwt5B2+66NaC7u0QQtoY+EkRB4ScamkBC5XO4ZQO1uUoFA292rnX892HyFvhV1e
CnjGr68YfXpNRQ91ftfbNNmZPFOpKQK3bBpsCzLka4wOGLEXx9xdUwSJBS8JA6DuOtSTQPyNCwwu
2QeY5ljA0nCW5GcS1uM/UeY/dRJ+xNHeI/Cqcmeuh6+DlK1PJ9/s3P9t5F8MAZyBqjBHvREfv7I/
4cHcLDnZ9looPKl7+oF5S5oyygLUmzOPgZagm/CuRpw706SOO7BrLjIIV+5Mf+65+7CY0+lk9qcs
m2gNIxw6liq8svYWzBer1TQ2nOpvN89gE5aNsVI86fxmrRGQPv8FyUS1Jqr1vcy3ZIQxB2qauuc2
8zR2LHCtSVZ6aEvVAUwqEQTep8bUD4aAt0xtl42hw4Oz3VupzLpwZbFBm5CBRcJnkluVztabHAFJ
brCRtQpz63VmsEsL0YlkeyyP7lntkHpTSlKHWoDsbWbm2En17aPZc2Zd/w8hKB8ZBHkDjbkhtIVQ
KGI0BJh9gp1WNr+zgkdbrZTo16ZDUfGd7KwWqNPkgzSykGyx4gvcVD313m8WAyP1lqBPmzMy1maT
pKm9D7Ug/ZXPkjwacp1KdS8d6rqwVc+Lu5wXliIKfE8OolsOyM3dXhA2Nc0cQ476BwIRGeNngUYu
5Xk5SSwOg/+Bv3yVUecZvqG7x0tJQGBHAO/9rxsgG4ebVpSI9UnQVjGzS9VNKIta0KLEEEnj/O2m
lB8W90eowUROFI9Q/t1Z3ZDsw/uxbV4hhyVLhMaLBHjwdy/tpeHW99vYvJYscZS91Opyl0pxbWnm
ZK+W+qBF6p99O+ruoh/7njGgpw3ktT2PWd+uaCFseZgkoE2FCHhk7Qsnx+jmmynVukKaFDZkGmLS
54kG+37bSfIBnwb0M+b2h2dIWcLwFI4gbOlnKiE5b3MhKD4hoPJ8v6rSZVYvOHmnkZai+RbybEWI
FAqhWdu5ovVtPtJGGfSBhgpT+vhvWiYbhgCIt+sxKoDdm0UQRrEuedrRHU2W6oDz3jWHz5e7iciz
DI+aLBUz3O+hyyJSINovUcWePlacOkI7sd5XOn5UlotSlCamAQ1xpECcSeWMJLPxhdLRqkAsP56u
+90CrrJda4KyY1fK007H9cUpyrg31Vpfwyvt9+/ncWv7PGQ1t/nhIHhP92Y/t5gNZbRP8oK3b/c6
qjfKfxwtTcvJStZUazSs6BVr66ULjNoKIwdxWohCRHw0M1k4k/X16mMdgXuotE58ND2jH1Y/Pc6/
kwnuWJ5Gd50s17ThDm2GukTkaaK3Kb11hmiCeUd9oaMeXdyXjKGO4Fm2NEmZOEv5oNgBhgyHKyxF
nF997ngBkxB0celsGMuWVTuBJROf6QE50BYG1CNgpUMuLnVGFWVRRAn4a59DAG/kiP0gWMVoxBVp
5MgfZT/lXyiJnslJQ6mA4KokxbhnMgmx5z+OY40UHlzlfyO6F5DKZ1/BzMJCN0f/LYod4ufKqpIe
DV1eMS/V0M7rAZf3nCwbIaD4cMyWUCfaBbnacf1FM2CbDBA6P/weqPRW7G1akxqkBtWVeIoHrRvg
TYrN2jwh85a/tn8F2d4Ku7dsBtA//UAGcY/OkcLV4mMYEa48ZfXUCEOGtsrLhEpqSwElj2zhN/zo
ucVSJ3KCTGaFOJj9UbyDOsMzAnDvQmX/g9ycHCe1OkF+hI4xPhwCWXHddL6UKfClHdo5P8RBndyG
cBW+iKkWWukOeklL6ig5g2jX0ZyQP6E1i+9WT3YBE7VmNmMoLLTajpNg5dCXsGwiUJ1ASPzKIQ4e
1jdPcme4qTQ+8VY67CLgO0PmeFJ1MCXvfkJ5f3OBAGRNnY5VgygYX78x5CFc6wqtDIRCcF/cj+zh
kcIaJK3D9YkkjdYTeMI1LE1elrwY59wzqt/izbzDITlD7V58nt6clysfgoxzlDpH/gzx5aJdH2tE
8hHMeCfAW2QHlHxIJ+NQhMP+NxZi+EZ3UdKmfvkcIPhI4pr9dNgw4B9BumU1FRA40r3ByfBPb4/3
5vonYs3lIV6eIHgsppyWdrkdksNb4UrXhmJI5HaOq6q0Dtgs32E8laM6B57oNU1ia6OA/OvSVef1
fy015sdZgpu2sBiOC6V28QzPHfXIvh7M3+Oqpfvg2eyOkFEoYl+d8hGOA2HcCnc69NydWVua7OF7
DTzDhF19ku6x6DLhGUUeEN1Qy4Ii6NFJY+GqMb6hIl0tLmBa4CBiVSIKvnyIEd3S0X4LXXOzOrqy
89lLSuNm1Ksh9C+7+gkUzEMmk0/l+xfSKR6ioKslFOU6fXczORdMjIRkWwDhqrcbrZVYz9tjVhn9
OKNrRDfT04uGpdsW4vSiGsHj34dqo1+DMlqL+d1JCY9mYQfPCsDYJeeLneztXhEnnJrA4KGxAcqO
44fmglVdz9Zzll/ccjCPfPGdROQEMXjzP1zbIeNsLSVj0EqDzYEDjOD+AsGpvbGIHa6MtvbS5DT8
H644BXtAjKjh6rPAOca1cYMNW0QihAy1JicyXHT8By6mxTAaGrJGkwA00bRVaBZVMp73oXpYDkyN
Mv/jRUhn9moShT11Kv4c5s9IVfy2Jyz4EoUquivhsyFmj9k4eVNIjOOmcPQtB62O+2Gpts57CmSC
oDoaUZf5qEQEK2lopaBkuIjabdx213temTBB83H3os3/t3twjbdfPQVmMkM4wxpjOuX5lJyriq0w
hUWjOG5rAjXBwxmBYfZKvd24zznCD342MVbnsLlm6o0Jrjm+0pwJjGShKMS2nb2ntZwzKlYxWzVH
X5UHeZYph+TFdf1s6bCvbHlpSvyA+z4e7kjKddqdesLaQ7arBg4Xqppv9HpCcIRyDeJqPzXfP5n0
OwtPt2wYttUzojUqF+ztTYnjBbMyK24XzUmix8xutigCV7YN5QaoZjjaDV1EiWbbNLuLtFsuV3sd
iXTJEPBvjGSsXQDbEjU0awQ7aXclJQHog/ghSgJG8YQgnGyGl4h0UcnJmgz5zlzCrO6LSj4Q1VvP
c/GoB217ewdNIW324CXbqqdpdvfbat4gZOUelrjVVUrqcaiXiCTNI8/8ThWUaUAGCo+kdNbA/+Vk
xrWGZilqQ2klevzQbbVcPe/K+/wvJTWRdr8oFX3cR7QygxB51PMY64sPDqTdiSgkKQu5LyTTwBbz
SyEWxZlp7ekHl9svxGxeFBnv1LQeJn66tjk0Pk7YPx1VyAm/zkhAGchLfF07qTvdGr+TdpuFGdhb
LKpV2dKrHxL2qhlGkbj9XP5SJwNmJwwmDv2bI7mwOwcp6XVgPMr2y4Exlo7A0cTQ4yssuiSZoSXo
6UJ33iSGCxSVwMSfvaxkMmxpqOuwOJoBa2Z8H+B58hEfHGuaVd5gkC78dlr8fgjZ4olI5rWIbZYS
pD6InBJ9YrMd/Q/jfW9cBkmJQkCIGUnBfAPCmYHGT3opvrJLI6a6/k33VJ5yQGSKes2x1Sjn7oU0
MX2F5zZV+hQHzy++JPo4ST05wHojAT4B3uum/0F9m6frWiQ67Z6hI+Ftp2XOC6Z6CmXxwwPLo9tW
20rpNobQEQDuz9SlN8C5lEj8e/LJbD5eFc3fExg1GxK5/Wg+KDs2Bi1vxWwlpILcIub69UiDz32t
qPdBTpCzIy4a4tJ7CqhwnvUnFjF0t62nselHiwzKTkOqi2ezi2jZQ2bR49gtwbo9PNJ8IzoVJwOd
V5OopLVIXgp/vPRJg5pz2Iqd0fqtB6UdLQJx4WDxTKPk0lB9IAXjuBVepmzesFKRhyxOXTgLk6Lg
6EyHOpgUqPqIdvcGYLWvAslAlRjeoXU2tCfqTj8R+iIxJ4qnu3eJxGV79A0SE9Wemi21/FACDr22
ZEzDTeL+c8hkCsQGiuVvt2sSQ96D3OxSCBlF+MTVwjG4fa74i+60wdmcDeYYh7wqRiaTOMiOjaY4
dERF+itbkVQt/P00kXJ8Iyw0bkdzSqu976V+e2q8zRwAutVy+Z6WI+2Z4ONvG8SqeTCJtjI11Wif
XtBYUcFlgtYOt4J8M6v9Qh+W5Xwb0UmZjJcQJTmOyTW3d/yfnR+uYF6VACM8o6TDvf34zGncaX1b
zaNRIDE9K2wR8Q1APlJAdXZ2JNflnbrcqUwRh7WoTMm0pGwMX0H5ZRkVncyLIBkzhMRu6X6AkUSg
BTIgXE1jZebOaZXdg3t6aduGolYd9rRFpNtKUgpNzEQA1UZHHTAGNWK6KHo2DozUdZj5uGvyqSn5
UVIAiJkSAyTbcjjwKoGiJY2kfkXm18fQdzCwG94jl3oEH60lk7RuKLVPpm77W12s9pHubOGWKTyt
bDx/cAqbycEVRo6fzg1Xrs5FezVaRfrAYx6mBFx6IkGE9AV6IK1B3nXTD5bPGfjPJmZhQ//SK8DZ
/SY4/JhF7g+VynA0zydQQcDXsXqvHO01m+gVfTVnOc4Wsk13gEK1qb1aVR/O3o2oIs5EI9vinjlz
VUhemDvgoOdR6aILu8aW5ebVpnnedfdHzW858bDGqejhp99/epz0/AEQNCewKGpqH/LS1iduAvvG
wGGgf7f0YzpMQIFK6SU9T8aMBfr0ZO+/Di8/Jwnkx1xZn6Lt7Fq5KIc1bVGjoDDueQHVpdM8GghV
b+u3cjgXkyDQeR/pDFCNluVAuDsbWS2pWK2ZLBK27e9MevBOifWMavStyUxkncOEd0EsZ9zcGvVs
MZLDGKzjHPfadYbJQOxigvybT5FajXOIXJPT0lEJ2YhoWSWeHJMh1ELfZXvJ95h3IfoL09v436l1
d15elzJTTwC9lKOJpTywI9CzKDR6ye6AYZIIRPFb73xCsQqN+8SdGtF+0YEaWuzQD2uEMtOb9IMi
DjXJmu2Zbe0imGHnwJa+T8w7SRjeWih7WpVmLVjPjMHEeIISWb+lAn1BvLC7oM2JLq5OvR1UFMAN
lhTbw6Sf3N2VRVxVKgtmMrUJk16+f0R3Fpg5/lrc7jAQG1DGfaO1ododFutaK7iEQVxkXUOv9RCr
kCVB52aIomSJxqelPC811t/vJfR2KX060jMTud9bhECtVlqd+hRw3QmTAmhmx+1f/pUQGcewhU2i
OfqdBi6v4Qw3X+YkHPQ/QGyiAU2WliiER+NkeSHDfAsvw04QpNZUSy3Pae1P+W0sGLSalXvp9riR
twnJVt2dMXAYOOF0EYySSLlmD/xRBQ2MaiUE0EaSJiWJ9Tv94zIsDHrMIxxYc/C0HqEVC50Rnls3
ESt5/KmKUDJSu3Q4IhsMaFjABEsV+zsrnI8GptIHySPCU5mOuaZHhHdIrRCkegMd2IA2KV5Aumo1
Gz26vYqC2EXVIZCw/HJ8FMaUrUv+a2xOSbGGpJNeZHwRItWBQ1L+T84ILrUVjq4qCfcLLSwt/Ut8
FwNfUtzmCxEZyeM8CrPH85in3c/QQ/hs93yGmqRqUQPXaxLrUKjnL46yC6LMJi1Uk8Ef0CzddNxa
uxfZ+1FdY7BSYgRdCfDqfdiHm/u7V7DRyCDoBLbZSo5wAAjlWpIC/aBZGvaceE9xjPeUcy6Dystb
Ck9B5tXfDDvDifRkJC3eU8bX36lJ7xxL6HyTFg/AhgsMtQSa9CbIEo6RtQPQsAqmitsTzWcjzW4z
9JKI4L+tCOe5IHsZ8J3VdJG66CiMDpzaB8DN66RoCRm3IAHQLMkTXkB4eTkW7Ckipf/0mfQKFd1u
Ss1IuDL+lI02ieLh7opmB4sJek13ISw8P5Q8l5/x/ALShkDG+mqkmgZ6anYDiTF4n84GR32P0FCR
Fzr8H+H3ovvQWonU635btW5g/h0scWCcYYDmpf54zKwdSAekutvC8Ob4irEoZi6TreRVtvBFujuR
DvH+fDIYlHr7dwI/D3flw+4CWp7PRMztgOdiLac4ygPM7zaj0DEsS02LRU1SQ0cxRIV41NOPBXHj
BV0ZDEQWssGWWHcsNHgwmKktUDIGEFUt9DaUHuXAy61b64dVgykAz+vf1egvYgpruFlglpk8tj9T
73pQIPlrE+vC5MyOskUzF1x96e8y6bA7DVhHcfZiR9ai+1eeq7ePYwbh276MW0UXul1K9s9Fn4fM
GFhS5BzMxPB3XlnHdPLf+25ztM6VL1cnDgVgiMTgvg496gGSauX9qbi2KIz3hEFXY+NdRE0KqLxp
BpEvXDpUp4j7YyZxiXzTuOUUAwyIAP74ucvCPzW7+1D0nVUNvICZqO/EiGBXGEWzrojaazu80XQk
vRxqsa/vwtLCPmM9RLaXWVRvi7+XephcZzLIGnkKUOkfwE5RrLA8uUfDIs3Ry/cM6E1DpLYXOQbu
Em8Uj5E1ClkioMSHrr9FsZhiG/VNJ1Gwc4pq9neOA4nrBdGYt2nh8L0X61WYTsz8nEB+u+jcM4N6
OxNBFKuHc9ushT6g7ofxsIKdtTrWarM4ffzmom39KgEi1s+FB2X+K2MyYEpXrc0rrsqjxevDpvqj
0HPSXfuVcGif1Lfyc8p1gwubFNlIQmhLs+uSdFhzY/hI53dLp5Qcet6SORpPX9eElqT22UN1/jGG
GWSowOoiJvqBMCGW1KVClvNqIgsOFL4hqHF5vq6vGK4qMikWntRjp43mz5lkGAvr2ykwBU99AvB3
WDtQLs60PQqWb6lCD0SkqPuy3M7xIjIeXSIXS7Ul+SI72VW9mZkCPSyzzF2sZwKLC6kiNgWXQ352
6XEVE+qqzxe1EbntYXJLlNE3ApbbaXfBQfMxtlFuhn2CCNszuQihmF9+ql/fuEAqCX8MZmv/ZfIh
TvVymAujxQgq/v8Vidwe9gibmSnVQB1diYgoL8job6KgAUjjZsOJkb+1+X77+cmwQHp69qTDulX6
1LMAXaEHK8+9q7Om5NP/kTjImHwNIV8eez8+WyVpetr6kBv9U3zQe1IzMTZk8H5D88JhBb5TsIoH
yF1hd46DAY32m1w0h2fTQhPZarIUKRU4YB+s9e1hNzXykcSb6/U8aRJlVdpTJyY56+/HO+cC6y9z
b3tfYSkGHZLWdlkIGXA38cJauKbHOtnLJMGAYOczz7qR020VZ1XRE7vM/eAsF1l4CzRDyRtUNYAp
DWV93NmKjpO7N/B7h63LBwd6t0jvxFZiAsnMNybStI3UHgtaJs/gT3umX6J/XeijHpg+ACL0CXGu
mbItTveWWMcawq4BgoppF38USJOyeUSkjGmG4TNpjQzpjOTYgBwGVd52fNG3NeQAg3WxLuPZhGCF
lO45ITEMxjdM39jclC9hxqpFZ95gQGHHRILq7nlo2eW6UBggAB+aNyPAJL6NMpVzyJquYfN1KhNZ
map+EongqNPrDULQF+HWvgbOw/ea5fSrGeqo10jJcBZ+LgaSFK0G+4VdjSHVfdSuxHmJNX3Wwfes
0AeZbb5CJ5pstxEwX8hk0oQYd7xA1BRKMoAE8Mt4eastSQGUl6cI9PJ0rtsFCx54IfmQUdDQ+Hdv
4x9E5VwxjufY8H9hHLLc+d1i4qztILk3zTbz7kNI/HRsIB4EmND1CV1TEtchNV1RnIrtm82ppLd6
PtWqDqyWDnjyf+hutdo2m2PNOnWf/2msrhrEQqACmLwZwPlBz43ZJGsk4iM8/1LRPvL5h/55nS1p
YzVEw9HmyvRY2YFGdUfbfYWcYEvl5D4rmBaLP7IThFJTDVgHCBWIBmQ/yu0b0awmxafp6TXIqGB5
bycf9xtzGV5ugvLunVFoql8+oK3SYyy1xwzQmiK8vg2WEb6OvGp6FZ8mhPhYwIMu4GdnADwN9tGA
uhcBOYsVNOyR/B/V24dHGDwAGx1Z9+NHLMW7vd6q+w7NdYjc81Bv9CH99+bFRdUNl9Bj4C0ktliX
0VZ+qaT7xsttPSrusDvgbKEAGBMAhdfGikuadK6wAXPmLbICPGFKQee2/WvmS8r5rypIwRYKqHLz
bT21clOe9W9XBgvtGj0ql2sBtUwgwuxvM1O+kZGBlf1xVdOTyooe/3NOd9abR1YT+5/AhMMt79hG
QBoIRaCrIVx5+oP5ipAMXlnjBAwrTGq6lolUxv6UBKqQlUUM5YKkwBbTflSM0jNCECVT/YEQEZIr
XpPXFXDztTzKCmZ3zOBmNF8arrZ+ciW0EDsmxzOGzbmQa7fdjn6U6kqw6XEXPhlqLja+HGRQctlK
2lmHpOc0G1Ii0RBGHrnxyBuLmE641eeA5vNbpl5LPh5ZDZf5fOrOfQUw9bxwL2KtRnPOdY4s5GCs
mXlrPpKabSuV5ijggBzV0aU91bmfQiHu7qOLiT5bK3LcWZn5iiJQJ+W2Iyqr8/F0Phf/mOspAxe5
tCsK7IEmnNqonBhnyftO93peE3pOJmUP0DTinz5A+qgqDI2rNeXBRqkaugM5Z7yrhFX4ydZqp5ge
eHGT1PGa3zkNSHZdVc+SbgLkNI52DXBSs8SUGJAn4b306BzGNVj4Y8ZxkE1vLE2+8dqhDR+TnV2c
J3N5R/1tCNt4M5NzAbExoQ8QD7F3zfQtI4SYSX+2Wt/q/ze9tJVB0q71iYU9DcfcbywrlkYNxPq3
C0WoFZKfqaRdbM/WvkfARMf0XaG0V3Ywnflu7kaYjiHnF0wRtgY8ZLXcVLKdo/uE84Uv0386H59v
XuFaN2BoYE1QVa44P5eZuYJ+OQ32Vip5KJA5XWmLNy2ZnB0zucVHeSQfLuAxwRhsSqFFXtPevElB
zSlJ/zkVJFBTHRAIEg317SKcJ+T1GtaX9K3jCEKtIZNfmuckDOCmtUBD+4iQ6WTp83Jli5YtJdB0
pJfgIV+rLPxePqycmHBw4ky7dP3Z2N/A5PTJkuGlw1BkMgcV8Iw5NLcSgR5xeLhRz3IYjZO5DYSz
KrxUZXXRb3kQGFH/7bOdTfXB842z9lA9r2GA+5NvgY54Yb6McahptOxNC7Kza/08T4qlsdqUHsU+
ZxX7XX4+LEM15HSZvThc9R77LEnViNDtxUfQnWDHbfYBBljx6A1OoFJ/3w1uvAr5060fDUacoNYc
olvHp5sYLutRXxvhsaaE3xSrZ2Jj5xlIof0VO5W9CSG0ZYpVvhtJzs+b1F7wt5OvmYVsd99OaM4V
BYhJrTO1QGf/XNeGJxYRcjGBEIsOecKNz5La69GL40O2ltdUmPeFz7eI2p9G0jI8vjUF7EgfZMl7
lZJRBbk2y1/rGhmBsY/810sO5hTNLjJcFgvmfNSgRRJ8bNuolf1qMMa0WcNPahRTwv6bxheMqbEJ
j8T39rs1NAjhmbQZgfgzQZa6pHTh/DWTab76M92SbNfugYBruHlXTTgwiqToRIh7gdirFJXXTSCC
dtZa2byMGCE5UeECHM9AmpUZpFMvoyA8CC8aP8cHXnjNebW7SJvQEVqMTRL05eZAgdhfl8fztdeG
zAHUEnjedjrqOl53hAmLw7oln6sNnw/8FWuMLi74aXjlf4rBfpWmnlzBPe+wT7Nv+a7gcGVRD35U
Km43scyy5Zle+YRQlkH4cZWFNVTXR0xLq4+4ZKWeY9k8fYcJnTmF3b5I5NzG670bVoWcM72NGM/u
06MPWOIxyo4ET2dZLcBuC2ip/gWnIKi0qGFp4EiFkdjjZoFdevOvuG1X3/3epcyekkaf9Ofrl6+6
5Y8w+7+SkAaucnbLOSgtO5DldKBgcHMQqs7tRPBr+xOsB0pNUCcIiyaPK3QMMIK1sV8bO19tWYYH
cECNrC1AdKBR2Ti1INesw4loghNnKbrEH6WSErS8+zNFjoykX5Q4ioPoi1jdqeUvU61TSgkC9ptV
zEKYdabDWTJ61h18hogwZjoMMpx9h7JhafpyDhm2Mej3R8uaAYIIWyXiwABLaW8sMKjF+/RWwa4A
y4P6dq5MvwMZHpRId8kj32xEDjlWTVHdY1G2jFN+uKc9KjsjxkF0s6tObFqskvDeUxEWulackyea
xIf2/3gPQeVKIt8RHcjyzpEhJcsIcy+y99KFDGJiwhL95XpkMBgYuKOcyzcNgELnm+5IYPKalm3a
jASoErECmcwqWdLWX81buRIrR/9VFR5qbWAmJe9NgaB8RorrtfTfKOqIebLuECblixKrMDde8dnU
GIPtqxsVCSrk3IfAQGoPdySVoGt0oaME/tAO4uK49H1b8EI7FY6+vSGsk8/ZNjwCKPqrf5NjtJ5a
itElUKNd0XmUgGI/qngl/cpncuXIkEcnvR5DQ+ZERY0w9J9rX8ABZGae704wwRxClqs7jj44FmG3
ZHrWurWSiECAZFEZbsPrS6mwlGWwsW3wxSrwM00rZxWfg7utEFvMhetF/BUs0J7EiKQjj69UksH5
Dhg+jqnAgpBFSn4kGb9uFR/tBcbnVZy3XYUD/UfN8G4s3sy+w1t+Q5dqp/9oRgZOEXhmjdUIWG8A
Lezr7rUygIVrvH0Xe/JEdrabRenKs6nl6DRuugFCrafDQ1JjnHQKHMziPdo0XNBMc3w7FTm+FU8P
DF501UEPXqWc/14Mb05rQcAKnOnoNLFbspUTm3PLPX5z4OEi89FIIZPHKYn63gMIQ9EXkvvBNJ37
yaHDM1Z8WfnYf3874eyLXqBC6olDF+wi2dR69gPk6VC1FPNezOmlrbvJvLJxDS/wlNMGiipJMr/y
yiAdVW+FG8po04UjKCIxbitNoHb9jYTEUNb1Lccw7MZYKaeyCO2J/NR2zr4t0PAtZMNNgm/GOi/e
6V2LVrnmlnLuV1EK+BRBxjaKgaRrH9s/jzHQfO+5yhVlo0Q5G+Tg/WW+qG9oCqcucf3JNoXj3Jii
ekvpWk+QRUfG4jH6c4TVI0d3/3bfEcwC3O4N5H2kcBc4koPJ9igaIGsyGvaYKQO+oTjSlBFz3WSV
Ize4MkAP7xnI7F5KwSvLSTCXHtRFHSb1M8UNcUtlBtPWkyi6sU8fvXfC6AlP4Lvfoxfx+RHTbH1r
t7fnJk7x909SKkB6tO30cl4ZC7c+YwLTrHruI2nr3xAjwx5mr1nMYuqxRDFOrlUuzJx+ER0OH/ZY
swFso7wo3JkYkmuZtOU0SYen8DhetH20ts3HAgDcvP6r1bIDZkNZCGO8it+sKjqiWHDkfJkjXw28
8L5gGvG0NZdwmBtJI9X+lVu2EymjwUVW5yb3To1CCG1VdTYDZSh4OWVb2ir4Onj0Am0bVGd+Fdo2
n7s2T+f8P2272hC8cNuLeeerpu9pAeoCWuKMGBSEQJhLABz01xMR4jNLknQ08F5IllfZCeYFGJk4
My461jxsV2fMoSJ6d8ZmUn0A1wPmpWL7c1XgR4mO36vG03V0BKqGDbOc0MafkPyPe0hk+BI1rBP5
mZz+FrN53PxC1nT2lWSjrGU+cawnk3ENUwAtyJJ1MxVYbCGQACgy9njctBuVXJksit4w4PgItLT7
yWvj2zVhhHQ3vIKKPiMxvGQBoBgP+SUNA4jTaa+34se/BCx0Qt0cpkrx9dKHNqzoxJWY2RBSwdEf
Uca1/AidGWttjtbwSxCxXF1BQwoaGzRF/3tf6qiJmjp6Ptr8GOwtGiB+D2Xb1HoGuR9fQPhb8Y1Q
EYmHZS+xVRQO/c+zPBuxwPx2OfU9gZZ5i0gMr7y1+cwGxnKiL1VYp/epF8c8JTHBnOvBEA1Iace9
RLT5kId0dbk16QZt4CcYmlsUK8EG42Yyo7S5aRR8gjIUx+5O5OZmtym5PBRmHQ8EPwdOxH+COTz2
vrCdmXxDjXZQ6vdHv9ewMZuktzggbrA+84wAL4JdEQhVaNziqf8RscqM3fTTeuBF6biiwhWSEU+U
SQzZYl/Q+bGdnNQVcuYwklLx+q9hk+TjBZIuonS/ijcFV+1MzCALNaAFrl9b32jjIONRtsudxgva
gv3GJVTu1vYnRug85OfbC8h4k5kBpo7g6t1upRwWPffea0q6ATetNjue+GWE25JcFj+UqOc/+bK2
yQyh7O8P25DFq9s/qkXZEB0rJhaI8J4OA3KlbUYNNrI7S8GxmYoLynQ1wjGWl74e679DAIDTSkFE
XByjsPO2KUGaR54LeHeof6VLiN2JRE/AfvCP1CCp9By0oVMUKLt6hi3Cj9vqCVwUh7Fz3/uUN4ey
odOxQQDF+79nORRYNuiDfqN/G/AK7bW9oH5EKV6z+9rxqaM7jjDnl6ZTLadKCxXDRtxV6I0Ztrrg
Ay/R4SEfWo0XpRbT8FjXzGRqr9pOZ592ToN7AGiL54VjgkT0mRHp52jkBnIqYzYCNpkRUlz5OwVs
dpHkkQx5absZarMH8lo9WaAi8z2HiXOahSxT/9ZQNfYv9oZwNfx9kPqtJgWzFjyZh+0q2dJw+Bth
2MZBtEO3SOrnO7IP7FU/37f2a+kbSWIIKywekZRs4wYf7ru2hfFbS5aubx15U0lvU8GMhaHQjQXk
LpQyS1xNxFTWvArSdIlgOnfemRqM10WX0wKB5JXZ3hj5O9ScFTEs7rxvqkkVX9XYp7AY1tMeuiAL
Lv2uUIp0vJRsZ9hBxCOzIC+xb3LcBgNDGFXF+CZSa+tpU9C2dMNKxDqKy762EHu0p17rwZJsI5kY
mqoE+GO7TOaMejBMbreJ/aOrhdcGg7s83Kp2eYMB85qQgAaCewDM8S+oPGNmnTHF5dKqRqRQm8bc
W5EOl0J1n+KXyBcFsuPdpGI6upZwEOpnzYlmtvZdbdSKhaAOiSQ1CZSskJa8grq4ICJ5gUqHUlxR
5tJf5mX/X0Iz5hkMSLMaTWXv0MA/UmXPY2Y48jde364pL6iztf3c/ZVT4G9BOW9WYEBYg/S+n7t1
PAezhsYp/cnWs4fpvMyik9fojkl5vMLtFtWnujmljCH+WVrYcTgn9Wn5DYwqTPF4yKf6CMy2rfIR
QNSr5laKXmbMWkIlxA8zs/1eP3vljybeUURNkjKz2vI0A9OyewWNOW82K81F/R1bKYyfLzMAx9fH
kvDZ/fQSP1Xv5nYBSvFCn8aon2IAcz+GzFB837socb5aSlX6ldtut77KhBZEg8v9Xqdx6mbS16c5
qSqBEluIlcPfyh8VC45w03mtmzYBtzlPDUyr7S5xzc0iHWnJk3GlDNqkRd7MGK9yoE3sjjMBlSgB
g0daL9sxULBRyxCcgCbLtNPDrgyF31vZ2k8BFBhjG4XA29rm9prgM7J/u4FTxVN9RlJcJGC4HxZo
9M0xMcnughkVCFM75iFq9300Gm8aYbiMAV9vjFDjL2wxa+SM6NA91qgI7yMwJrUF8BAUQAFRk1Ya
VNWmhER5TpGf3LSOhNXsYG00lmFvLceBFoGcWvNjpeEsn3QjNt2l0jcz4GX3BoX4gXtBIIOJmeXS
phjKHAeHpYOiwMCM98riUrNMGJahlZeArDN9Tjmdz05ulVKDSqwgLq7v3H7F5HhLERY3+P6Lk1P2
8hNHiDDdA6/dQ4oBl3IBlq7+tZLbs2ALBVR7QChD0Vwg4lIpE9uZTWvR64crGCxaqZNzZ0Dn+dgB
uhWegQu0hZXFjjP9vmEZC4WWeOLh1HUEYFqfCzNewXoCNuYPwcyJcFG/RAuhznUmGyV++USgWtu8
STNXrqRgaGRjKVISEH1H/4QwKRiyVL+JD97dW9mSjOjQZAli0CHY7wDpMqZ9bQ8v/D3QHIn3gaRy
FqswWzTHwI8ZO9tRB0ROzeRnEQ6Lm3dVIMS9AwT+OunQ/qQRnR0Rg/9Fo4wpW0sTYpZzlalwwtI9
wJhP0n2WaD0sSFFA/j+R+PXFlboxwrzhGgUSg73QfaSPhRQXr+TmIUsn+9bUrroAEAajP62GFR1i
GbRn1PET4o/sYAyzPtuTMBTygf/gE1w/0h/DkJH9wHIs3gSHuKU7NTN9ZQnk9caTySqRJb/4TEmp
zmIC93Vd2GdpfogmNOuQaM61sod3n+tMm1wf544QuLKaJBiyQMhgvvcEPEV5uxhhzwgVgwZhQVgW
IdR+87gyEJc0RIXwhz+u/9W1wBfTVaxYwBcCouKbrsr5KV0rG+rT8T4hhcQWFPHDVuh1dM9rO+ZG
tYBnAUJQ7Mcf0lcw3f7j03BwRnJkGaAkLvsVGp8WKTsAANX0hPxPYq/Nkwbjd3QCWK+w8FllqO9w
1vIbFcXPyQBSx8ZnoMPGL3ctzZ4hKMqVy2m59SNOX6fOmMKY6a8q4KajjL4IjAeJ8ngeHr/y8c3I
eFb1v+2Ud8Z0Wm7nrJu8el8QNNb4RPCIeYLCDw5N4H7Blod8pABRoKhZdHRUx+LXMGUSLKsdC7sY
r+RZWmDF33x2lcmnmxFUKVE7kCJlolx2yKKevrO/FHJ4+WEAaYxDa/9S9ahOJEPHd1WY0e0PUELq
HCeNLKilup4Toqfx1At+7gVutnEbSICiGkSe1FWVRWIwIr17M7MceuXj1fiME6NiDWJV40dP2Jmw
DiXwP/Rf77tFUPmSlWuS5RzyBEpZs37wdMs87DqYBeWeLbF9jj+3LH0ix1GjH444E0v95vN7m9Lg
8eRis+Ok4XKhr8Z2L8bZ8tj4VGhMDXKpsaoSw27wEv48MzdGp0eKhl6mvOu6TLYTgsYCi8hlpWGA
4fpAK0OAOczeDF1iqD0GxtCNZbH2T21ZBjuWJ8tp/gdHphK1aXtly0lf+4Fa+fmqvbOBOeg13BNh
8VinP+GqWZ6YTXxUhoyTwS0v5uN206fjQBXw/WSKqXXaiSTgvMmt89MaW2Ok49yjql28ZSnEFlI9
XTFXflhQPBGkqKaezrtS8OvodsBq9MDxuorwzLq+2nhXipKhFVKMSsCEFlhLe6fyXT0UCUUVdmq/
YgehRSsaztFK1658bJXCUQcG6F0E+zoZneUGENkGSTBHm2Ce1A4RMdjeyEvxxLWMtMkSVzyFFITK
3vhe+KRR4nrKQcaPmfOFlaYvQ6rNVC0uunRRhx7l8mniCBdD7u2W5Pb64XAnAIEx5aU1EmokCIUR
lc/rKkcEJd4TSlyGCyEdhzw9yYLBaiKqxOntisyswLPs/hyxNSNVi9Fhz0aFoRtU+x/gsBaGPfxR
9JDQTGnhTc3XQHp5fdK+X7gQvFYJeCAYEfvC5j2ugLrtfAaRe3ZdDpcU4uazDybqI4HAlcA7Mjew
n0q1uIpyi4siNZuN6Gbi43O6wYxq5Xkde+lM18aiKh/dvNUru1ZDOMaRs+7T7GORyfbk9gMMN5IR
vNm7SdCupq6k/GpyxhRF1hCRfEbK8i4Jm2bI8MTV8i5WguqAS/i6HIzwjGKcdDPcIIb57naBTZE4
BzSJi8Wh7+uOtV9RHx1WcAhyFpO3CV9inIQX0Vk2sdJUxOuXs8+/rSNqC4pUwV3dNhtdStzK63CY
z8v2ws5+sh5070EtQ101iJayXz82uWyhc2aUvcjjB3BLCJWL0itEjowkQbDdACMCKnpecQnG033F
YTdeRcfw/Dvh6VdF4qKccEcLoaHoeDw5wUz7GG0UMJESkpnLq/q25DGDW0W3mblMNymmd9xxZQUl
tEYuoAtkzxhgTTpbSaPFdb8RGP9PPxZ73Kb4vEWBFSi2K15EpZfK/+Gqmgz6UjCtNTLbIZKZJ47E
yTq5Xg5dUO8qrYOP4buMz6YdjYzbtUsRfFgwxMFdBryQQ3j34SKg9nxdf4DOUve9QGmh148Rqcw4
VSrHvaduxHKGELavcNls23wEiMc35MXugfJQprIdttsHGtT9TEpjlyM4+UHXDzgVI+V5Iw0CQM34
aMj+q+qnW1oVgzzR54bPK1cp2V3yKYIyTanUXXS9jGcfmgPHAh6PIj7aujCmowCV1gIxVDXT7nLg
UEbAaX8R4w49yzDHXjdYt/AioZ4U9TRfdb0rjDPmCaRZv9/3ehA3WZarkueFKCulsspiUmVFc4k6
0abnPNpGMGRWmhkv94GNO2PnTm8sI+a02EhckhqRTWGFBVXh6UAbZA8vJrAFLEfFE7Kp0mhFB9ti
eq0GrIY0Wa4UhIBJPIEN3lk9DWR8BgRazTH7ciukIMPl2qTxYkG47aUK5zaQ8mIK1ZLNfvBJouUM
Dm1SG0kQijZOXX6HZdsRSEPvw/9V7S0tuGzUXr4UE7LwxysDJMblQnp3gksFuCVJpgrvTbPdc8SE
07ud+6V3MuEfuvpcVTd1Owq1ibIg7hxmypTUJDCgJDn+WQkdt/CB8aFFBGIyaZ37laQbCP+he13q
NGNfSIEI9s9F109vCcbjdZcy7XAKKkz4ayhjxITXF7JmwIlolzexZzjoZOdcaQQjdoOjd9W31j5R
2DdZKMVx7XF72qKryYEwBwTjMOrOVuSaRjm8rdKw2IKBsL8Zs/DKKLFEvsC6JLjYCHNx+m1YnFMm
skoWDmoMlGTmcXzUP+/EugZnk8JPRELvCaOzINZ9XjvuM26Fdiq9P/ZIqu78LrlbOc1bYRAnL3sd
Gc4r1CSwFLlpceH8wyceeXKGWzrMVnFvKU9CsT0WCfcBew6Wt+gSKIM8K49tqv+gC6H4I91n8T6q
vkzmZCrA0R+wybxdperlo410MrDlM6prjl6wSlV65GcrxFWDctqIh7aycIUhjqZNMEZRU2yKLUz9
4LafslB8Io/xNED1UR7FuimdUfmM6EgUEM0ZJHPQGv9MV88LPU7oxVSJpr0SgbkjODno4ud9J/xb
Q00rG4YHzd0ORRtPxa46rXoJLjP6aTDhqGkMxnpvoE3UzzslpK7tGMbGvbygT+y9GMTmYpkeNMJK
WR/hw9NJV3XfXFfv3B057A+bfZGvbuQ5eDflY9eY/R5vHAjEulvQanCQ1707K7B+Awm3UIKCmjLm
IKhOKplpqpXozjbJDtYHp3mddaBTBSkxkArVjgEXxJEs5nE80T8r7jl4+bjBSusVmjRgU2Hsxrkb
uvI87FCzsP8xvVNt+7K5l5KI6ub5xGSRaEQLGbDNpdIgc6ixrEpLFyaLMd8MJxi8Ubi2fZ+lExyd
5wilKxjzUc/LyplftckJ8kwIbyX2heuJDqfXfvMLyi1Mc4cRKkQz302gdLRrZ9KkObRSD6SVG0ng
0uayMwGIqj8O9z2Mv+rURw6r7hckr10T6o0AWww1LURzQbtxX213AgVPogvmh8aBPEFNoSPUHBAW
oC4hQeCUjXZuten5r7pa5fMr7oiVRj9VmsFE8ZsRD6zArVK/Mv3xzedGfXG94IY9CjHaO9d8fA8o
PBoEtTN7f3czeIpF7OMzJR0aelhBVtzAuwDpE3RZYgQvcShOEvSZgaJt4XLK/TDgBBVuw84tVriw
wSejxxufmJwKfuL9ZfgMrZTT1bAOvTiJjAxfK5saiNuh2uCwSj2XnLr1BisG1QIpQQ1t4NRfaMhi
fsJq0fgU2PvYjWQ8zuVr1mvS8zrr/oYnx/H6ZoN69hkmdFGsKHDJzvEK9xuPzT8YywfBdtUrpH6e
WILTP/kCNZ0d7KSfdboz3Cikzc6U9q7FJYLJLMgMi8xENE+LJakw+jwix0GUFn+jEx2ykDC3S1pD
FCSCNQV3bkMsUVTBe9QSXRfUwhtLn6GYrLHBjhY/LZMxLSfvNGQUUy7OIktWMLsqttlCN2QpQ7zI
Hk2aL37IhY9i+mj8v33vxka4PLqjBx8InxtzU/+i/bvF4Fv2Zrqn+3FU5l94C1AOWG5hNBE5UxjA
4EA2d3NW4HhLrxwm6qoB/kfcgvySEgd83LFjYAQ8wpWHGEKKC/Zn2A0YYKn/peNhOO56bLgxDoSM
QnxrgVXHvOmh3NR8ZNMWnSHKMW8AoyCEbFCw67b0/zhDNb+3ZlOCO/z/zdJnHrx4qh4LcpYhJKWd
1g9x9foresIKaKLXPfZYYcYbxpWBPk4csi1SmjUfw6c/S9HdtlqLxoOsWkogtltx4IVt7oAgvRxI
a/Cuc18JinqM7BGd5JvJfeLVCobA44C7JS4GvqFPGy50hfm2xS1B7NzuE7tBZeLsMFEvKjHP+CMS
d9+5/+2tnzmoWs1qWPYfD1Opdr3LLMIjr5lIu4Bta5O/8q/Sl4kBj1902E1pKlMnga5OzIe9WPZV
0wNeseIr8Qcr/4tSjykdGMgUzlvvXRWwBR0rLlTQ7DugCGXYS2iYmMEjJMB0EaChMD0kO5rojb/e
tUaAcVJHIJSgZ7RfG5/w5dKlF1ZGxe1DzByocgV37EU514g0Em8/B51aLhD+XfivUMb/Swiz2MwA
PT3g2QqBSAW0wLk59q8WaQ+HmZlmtaHKMCB8atDXRpOiAEk0XukAmcE7im9k85A26xYp6BCXlqZo
RpeXIT9rAhWi5kkpunyWAbboBhzQ9fEzqirRscT+KulTv+/gN+SAnBWGI1541ro6NbNgGTc+XTLk
nA8U19F4HTNHBWJXQbAoKPGeLy3Uaa4R6RsH/2JxQy58+lEw70sP9e9QeaO3d1oMSpEznh/PHYK5
SSGrJF/M/+1VG5ZiNNTONAW1IQ2rg4bvTh5TB9IDVy3EZAgtHXG0eduHTqOxvWDEqtMVu5E3Y7jk
yH6u9mMcWEjbC0TxlQT7uCkrNpEb6V30di0LipRCS1FiIKhJSTl/2og8ZWIaKIYiSkAQ+4hAHMCC
HlwB3nosd8PJjkCYPNrs0NPjHFLqN9gVcOqPOSzy91i1zs6NgBEaLjhQPrvuXrm+HzaUdNr8X/TX
+o9DasFIBoKU0mlN+nSmhrMM7tbFXDUDIYBbTMDw+n0nVrnhou3pEKqBQ1cGXBroHBAlX72NgwIZ
L0+M9Wk6BcO67ewoKxuHzL1OxIPeo5ANivE6AI3hgeop7H1DDGnu75dqK4h+U9m74BHP0G1fmXW7
X8KK/T1MyRaeZsd7APvOYsVKpxVn4shsIpan1ItgHp25YyyVIyOkzi0QdJVRch7lZKs7s8Y3nkpC
oyrfjS9bn84fhZzQOSWRfk73Ikb+seNNb3z/B+doK+YxiOsSizmVzqbH2NGG3OkJ8R/PLWHZy11A
uireWVZ3ojcyHztNt0UCc4K0UPxzEQtd9FwyvwsesV5ChDaFwT5Y62INLoXcDwtBxKazNR94A1pJ
O4k2jYV6WterIp/5b+2e/QqbWUfK1Iwuac/uUuHejxU0WLaveq+ClOcJH32SOUTYMZPajHzxpqQw
a7vkmTlMoMG6kR998H0Yp9+QS/HRSxMVFjzEwvQ7dA3o6ylbhsSoO2tt0hOboWGCyIqwL6Nkq54t
C6jR6y2QYRHM0H264LnqSAGYOKl0b7Nw5NYD7HX3mclY9KTg5zP3AyRekjG1V+AIaJjJ/UsN0+c9
9puQxs73ca7DtpS6zT6iZWflcboHfeAUUP5V5NqF3mP5thnFGQG8QSZAe6nGKT4qYR0OEfDEQLjn
Px1ZDU5w98ZF6h1rq9x6LtVI+EWF9Vgqi0QjDefikg65fvfqssUL2KjFqtitblpnAwr0XUrwcnio
ALSQb4nVqt4Iu0izLFn/Cca/e44gELxB98mC9KVe9ngAIURU8tIMH/uo3rT5AHv2wa/k3iptt28G
VRCILCOmdpdaokrL6qTCUz6t7mFQ/BONLu/2bXaQtZmiwZwt9ZuHMrsrxig+ea6K3tPidG3yxeBO
JLQ+AqarvNRu0gDSvhvrZz0iZdXSuGlByU0xTW7xT+DpxcFN6vcICQyuOE0+SPPcCMiUtCCuXhxZ
XZBugJdFZxhNIaL3zKjWQrVdD/CAwRAtiwXI+UHxZdBOOoRGGthdUYtTrChXW97BqlDaleCWWcT5
ZImAmf9XnyZp6Ko9uWJ5VdFDCmYsBp6CVU5kxdDozTCAT5Rj33gK5YA9gdZxlT24IRkwwUSLnBPw
cKyiaPQW/mCQXjpkC8CgDqJekyP0KSNXSczuTel3EVntSE4jXqj+jXiC4TPLtpoxqbRjSmUCfA96
qrXRvQm2S3UtjuAdcHcBlr0WkAwtSmX3MuXiTvpX6p7QkmvPS/ut4IwuR19YuTfGJuP7Txoh8vsG
OVd+14hiUks5wBCvsQnpDL735wcHQqbWTICVz8CqLed0Kw1oRo0wrT+cX/qAxcBubk67m6yLKg4K
ajNVfY15uJuO6AUBL3RdCiyZogEUkRcKooq9VtveayN6IUu5BkK0TliP5VCnYjYZ3pxp1vx2knXs
hzz+d4/xNPJBp1XFxXsDh4ndCS9ziuRlrakw4kt7qe1dagCRdaNzdff4xz/ncdAy+b3w3HAc0fuF
E8BhbgH5uEtdEtDjX8IP83wgJ8RKkMzaboLAcJW34jZF89o16GGLysQHuyHnBeRw7U5LXi4I+TjD
qSMxOqOJ+Rn4DohpUh6OgcyGj7jYCi895toAAEOg7H1aZKLgwY/uV4xLfECb2IptwN0h6R9a5ocE
ErjgGnjIXLFDzr2JizEtwxBtYggBX5i56HJ5A5H93tspsxUFd1qNV1/T1tRCOViFJVkK1xWaWZh0
DUxWS4iGXqeUXHnfKipO3YJs214M8ty3BqsJH4kuDDQBEQbcrd8C+BP4U+k9DHljArgPoBa+siLc
/81AAYOLYDzz+JgfQPJLHSWmpzwGHcs5Qm5eDu4EDytwCpNE/M8X9QZUF4aZAVpQEn/EulJcfcJq
jDjQDTmw5BnBoAr1OyhJZcNBRgoEfOiTonHNlbq08AEnRbVSvXcveNun3ciPrzKh937JGJhXpz6r
4kJW2yu7LsO/RBok0QeoUhO+E3IuDnNgq7yGcJ33WilxWhWmgHdQfZN6XPf3by4gwCO6e71dzZ4h
aHwyFRPhEzCGUUMBLY+c6BEzH+0FOh4t1GePw5g9glhCBraZlPUSuL5TxA8GVeuys9+uG75U24p/
vczpv6HJEzVbUnFCGFQI775gSoAL4NIxwEz8qvv2q0GADhjat/bjtp6154jHdQu/bliVlJxmSZCX
t9uYG/XJG/pSYBJT5ZU5+I3cIp7jouBcmr64Na2Nwriqc/4EopAR8YHSWOMZ429wbXUl6S4mdfJH
ybcjZ6w4MOBsqhrFOLgrHoog78n4R+ptlzTWdz6t7IC9KSyjDOqPfyvbEI4A+rsUJN9saAHPvhyJ
QLVFAl0GCPxQn+TighWAiWnR1IawTWwL4GMMd+C1JVu6KRHh5lFpEi+fw2m/bZHgtb7jRRIYjhMW
j6Im+RP2jPWZBJpopBGCWDk80iUubGhZzG7SxRp030ILQdhBr0v9AXHMuVKsaQMXIcF8hAuhlp4B
BOC1vuV1MD9ti8b4f68uhwBO7MvjIjy4ohqA2S8Y07ZS29fjzAowaXT0K3nFvf9q/cw4Qy3GzKxe
OjIUniuVZ5PzCD6rNb5Bc1NBtHOQWU5/j+Bitqxxa/WzErGq9USqlf9DULAyOwxeLXGHjsmeAUHA
rQ/TGhPF64ltbDeGVPE0sZd92hAqaAQYT1BaMu3+DjXMM26G4XDeGDQHR7EgPvfDUw0SHTY7URsH
hrHB4HAKGn6dvFRaCR4ywaG9UKrH/K0i9bsAP9aPn4UPqvFgiMeuX+oIWLkC6iq6ZBhxjgopseRw
+JHbSHSDlYUCTRUSvG7EzLiz/GFDudntm5aQPNrmYPj6gr7AguPl4ayaKk5jFIaiZA2KGOW2JawR
PNsTVNiIGX1Lu8RWo+fSgvtGoR8R8zrQaDF6OB3GgJzzG+EGhNwF6uLSuABtf0zfOpRbmyPS0fOH
MMrTqGErwym2XISLt0fDaSUPU+U+aMlEut/+qE+N6ubtIAtioDmPoOzx2gRKOjz7Divg9t5wS3OI
Ck4sfNZexO9d7FlP7qcpvj7xF939zxcqhSTJli567IuYjJysXhuZ42V3ViL332zPOfcJ9xNZ2eXG
guW+Jrvkb5fEaLPus0iWoUvI/dvIjvdDE1R1Q5h8XOrJEZDMIsP18iZCHwfYk3C2APPU+xnaK/UJ
k+qWvNKJw4jB7m12qj5Ap1TU9aMTlHl0qAvuGvmWWgDdAYVPPVaHEPnVaETQW4A990/8aRLkcqEB
AtsRSrErgEJJ8PiDgn1BwJMNr00v6PwxK7SIv5VGz/GG+PkxwGb7Y9MM4B5icaVyTpcb66vXnwdT
XsZkhmxXun0EyfyRYuMru+A7We3w9/fEuNjAQj2AQNU6hsOaUXAUzOFOCqF28+GlgcYkfBm16kai
JAj4AaO8QY0zEf4Yy15R3otZ42cFD4047Z4Soatne/uAQY3st2tkoOdvUo3dH29TvuPnTm1F4mcF
/a3C9Zn0AIXcBWDw2RL/wLObS+fv0qD9YPDyjKObagg4u7QxgkTDMvc6VceAD+1FZE3P7ZEdgntq
RNKqDk6QY2x799Y9MKaaAt0YCtQ8XHT9lyHeQa6NG+GvuhN9n2/rPmRhgZ50hdLWVbfspYwZul7G
xEFbWpMovRZzXShKGASlZfSHtrvT2IJfzd9lm7QxZpUpBBVJGPWB7IxlDhX8eSM3NLtfjYFzsMQG
tCDrcoo/7svP3TtIAaT2sM1N3OJmyo3v2TTT6AhptWpE/lXTl897yDhDo2vWFcnBrNVTfhf5YTLM
ABJ88idPL4j//dcwxunEi/yhXrNYNJmlCkaYxDwOhJ4a9BARGeDuKh9Ap5ViojwCn5Gg2fdcfYvQ
MUtHyr5iW37+w2AbnyC2qv095qqDn/SqxnGNgqNWSdLb+uKlRREqOPRTgYGRrnIhLdHjeyQHILvz
CO/liIixciEK/CPIWWK+NSltoShS5JvK5mfceo+69K/mQTE4QeQQK3MWCwzpZno69PVT/N+hmXk8
ebBTanvANtBoZPz/HRDiwfCx+IgtIsvuofWSAtxtwe99KpXg9i55UrRSccm7Is4bhY0L4VhD3p8+
9h+DXj9mWFPWCtQsxiYnzdLPkmID2OTY6Y7feG8IY7LUMf7C4n/m4xWDXIq9a9mnE2X2qPEYZNLs
g/QEF3jMp6+pu8jNKRcdecmOuM0P5e/8U6nrpnLEQS5KO2ZLSIlApQh7RjCQ6jzAe39qIPJOaujV
VSob1qni0CA7Mc4AnxZyWJ48ZixrFIOII6k4H07MR74GaG+/BlUse9HFvNM4Akgjj2U1mcShyv5K
3D13o0/jbc+soYFBKDooThik2TmqQ6KoNT0MUMx5QNHSekt53ZUv+BUkiIwVzMqmV11pHDQyqq/A
U2rMSb8qxdva4YTq4AH/UKaGZBfaqNxZdJcuQ4xaxUMvs7gDlwg8cXc1Or9DicqIVF5Ul4jQyAlv
bu5o0b9J4ZE7u7qOPD2zB6bA8D/NrqV8qLgvHhwRCuV6YgQpiZq9fMjgJJOvSBXYMG0FsABPAJZI
9b+NPLSg5nFK9H0v0XevnMUH0qBxUMEo6eQ/o7f+ewO5UlAqhg43Lst+m7Oh+CFakTboNiNv3NHB
EXQIVMg85zxnQUGBzZABQM7Gpg1HFQIdf78OyPZsLc1gax8pXuqFWewunUzClkeRm+12JKuLMkjB
6KDUVFRCqOI4QDp/z3qkP060RbdRhOAZseR/MzCmY9xqFzMJLy0uEDyZlph/5/bRFejochyzs2gB
HROC94rDVhOlvvtu5+xvyoDXGFcIS9DvMBGxx+IXI9bxL3WafGjZI4M72q1WuWpoX3kGvBZabiow
QPR3aAC+2czBlbD6PElo7rVidr1wO/5SX5o33OvYcFT0X6ERjhDSSj+EY+LtbhTvbMfONtXgWVKE
brEz/6Ple3ligkm8dSWQNExLhR/SRDwrmd8H1lsMZf5LXNaLslyBvVsQtOySJOureqJB6iRdOF2k
kZKuRbBXYuC/v9JAnO4cIo8f9FgvaGWE6Yf4m9SuSP/AgitTphF24waW9fz0rWU74eo1uQjSjmfC
LrX2YaYJz1dAYV23NxBcaSHQsOJu7Ez4UEbbiXw9krDEy6jCgyQ5TkevsH5Lzj8HrjVip2Gsj1Lp
HsY2BD89yasHSZvPTtxqwDtw1BQMUDTGl7msCz0931vb3PsRjwFS6mJiRGMdtbIFeg/3WNKMmBYV
QDjMbpIfiQEK9mEHutS7PbzDqFbzTDgTNMd+pMA5TlzA6gCyJ80Na7NaOOrrUJzwJMc7Bwoc7JXk
rqHiZw3EbaUgwu6dZsvHEZwAL7NbNURTSxyp5l605ZVW/NftYXituMyGI1N28BFdg/NTWVnhjtY/
g76Q4RSes5otgAtue8OOc84LAJIg8T57tUu4RYNtJnig9KyHXRrVUf1eC57WOua9mK5QSTLyDWV+
hfMEJOZsPhfFzGnLXKygjPADAybRsE8+bsb6ylJRJT6tP8jimf1TdKfhNbXDx53bEDXhPhq+7BiW
zx5gOb6g85nZFfZJO2hfeyNQ32XNouvLmpq6ncfFjlL0tJzJ1WwggwMoJbee00qvPLszEI6lunCD
84ybdxlEZ+7f+WyKEMNkeAYtqobD4b6IXGIHRERzGrAOTF3qxeLsovBshY19OLxc3acDpCRL+gKc
UWrZyYUPKHcwB1lKovexCZZ3DK4sfNOqnwyWAKNaVVUpPIcRjtAiA6wIlLOqaSccMIYUvJ545fPR
rPKe5kfWJGPrUOugW2jbsdoGeOExyxM//R4goFZ8spKR6urMAyRrsLWxCdJUi0xCkYMLRpVYy4j0
eEbjxLNjwwF3njAQc5zpukFZIsurMV9kN4yDjw0yG+/W4WIBWrCvbOei9DmhYRlMDqYFy9/7dqIE
gBrLVidktIwSCuEDKyGhlIz7L2ZihbOTilboRleK3GNRJGhrjFgfsPeMJowhndYyWyCqAvUbApVS
aGr8iM1UT3L2FgUAt3c8n+wb7s+7jIUUZlEBWdg9P85daKDo0JvaeQc8ORauZDR34IDyKl0qSeZZ
nGHal/4RekHQpD4ItAipbglhFKNyFLxTEf4tdprM7vC/2QQMfKgxQk0UuKmi//H3hgQeJA5XZ40l
ycNfjszblLspT3ACrqryW4QO04mD/t7mG9vV15qrX1lGn/ivQC3fgURi+6bVDIjwxY7kAvAvUPfi
Kfmy1q4RPGD7dR0sw1tP7+w0p6y+F8rDx9CqNNzXmwyvBIql6CUMoZ1M7UGgDddQZOULcCETQWW8
6mrlW/qcM6RjC19+LGHS/8072QiRnbGOa2ZCR/edhVnPbJqzRqyOOQh6rKhUJxuFESCa44QVKZAW
nIu3giGDKqVA1UKGO3mK7S/k7SoQbTn8vG1WVBwxwe+LFa5AMDZqfrGgFmm1FImv9XMzx2OdmQV9
Yd59SGoH09jVyQNO2bi95m0LIxL7w9aE6EnyT6E/mxW5tasnS8f1NmeefSJ5atuB81N1J/8IDP0i
/1o6YZOA+cXeySDggMBZBrjliZkDC9Ynexc/C2K7C5cMWlpQsbp50Afw9R73i9PsLVSwRzUxeoLH
IEKJ/vhQf3Z9B/Lu6B00TBNLW0Ykl3qQEoM+oM7OaOvg6F5CXtxmiIG+TwCH4AL9uBL5mCoIOqrY
fWynbw3lINldxcqZh6LbBbHIQv0Ke+FDRFwmK32W8wp5kbyxwer7TyoSijBtcYN0nRnQrYFVMgKq
Sz+pGu5eDjj0T47blAo/sk2EHFbDOo54XluNUN9NZi48BaHEOYr5vMJSa+oszXrXXCHcSwfhuFAG
MTJx/iqBRI4uXLs0IiRP52oj26Aty/q0W6Z1nl9fede7qt0tswnbmza4p7bjgzevf/1bXNDQnXIy
0dVNGT9uz3uWvwV43VX5v4dUFA9/37BhfhVo0tfVrV411l9YebbNYy1ygC1ZKZiDZPMkTR2w78SL
nRsWXChcogQqVcYCWY+YD5xS4ZDwCnT4g+6+UZ110Z+KnHqG7ixZJ3Xmn89Hxtvi0TGv/rRHHtcQ
AAhjNRLNablgz6jillcUqL18cgvKKyrkp/9c7QBmDYNeE9FdOOFd7xMYEL0sgW8joUg86qYJN+P6
7PUmiCj3hQ/ZsjZtLg3JEUI9jJtapc7JDpK9IZUzDY3E6UEtjOIRJSjwjEucbxRA0wR5+l4rj04i
H/66u9jvdg3IEil/Of2sp4DNu7gxpec/8F89RzyVo+xqVFzkF2ZBYebIru7KxDlkzVRb9FKkYR16
bkux1tfumH2IekqV/zCmXgprTBk4W4+IYjx3inaX/vbQjTmm2U42woAfVxWPavBp5629IaKJRoWV
vbF9HpIBMcBvk7C/dLocpqh9yqurHSphiUEfK63ZBDNd7ZVBBrzz2EeGZUy8Pd7xyEh3KriHI819
yJob9tzjufj2kKOaw3MlgYdyb/bA2aizxv5tu0gGvwXti34bEDKtZPvqtf1LRxacx82U4PsbrptQ
t1ido9F5z2OGqI9KfDFn01H2/FGYOCYq5Pd3YPJnDs0gFhoEPsQz4EOHDfn84Xc4cVPRHE9x0079
6VRZ0NIMYQY7EMZzXZsV0b45Z6RB9lBmd4fMOCcZjBW2bCYzF9aTl7GoET8YOhxqx6mfOMVxwNj6
FcsULfbXUGoahWDnL+6iekRR72+fradWPu7OdYzPA66+twdTNz2RkKnKo6s9l81JGx7SgFczgDxn
IoPqNJGSxd2mUyQYa5lFNqIZIK68vbPR7o4bUmwIbNlwkkeVzcx6GAIUz4Hk486PD1+vjJyw1IM8
JiAq+tKr7A+Zd9HoMX3dainN44UHkcq393TOWN3dSRepvqLSvLKLjMscGgOdRJddmZPHSMzBnB7a
Q87BwNexKWFYAomLhW2u5m6mwhTz46K71MMF/cB6nD9AGWXI7pBeUEMAViuH9x/NIIrvT6JlGWa0
H/p7JVFv727vnr7nOUhCnkvVPIuwlfa/2YF6Z/v/n1ZkYOoJFYGGKcVUHxWX2hOH31bkJSsr5zAk
vpsHDDzOSnDDzGU0SdL30m83UZ/VyXPzvsXVZ8wfYbE+a1K7HW9IQdLL7wGHZ66Km2x/9r+YJh3R
NqSMyu4SMz2U9t+971fjjmF61ilTy2Nw4T+oEGI6BlUkqF+Uix4BCpIz4DSjwZwtFIAVtnq3fgiI
XEVuCsDIepBnQAZPk2BQEllwWUGNHIHel/y2eCfwoEuCPYCs+58LXV/0ax0tHweY2rB5EtBMKu/Y
5qlkYD3ZRfjOMVSm8AhZ1ZomPrXdHsYDo+lMRwzIlOIUA4aEpZUWxV5ZfPA9/2k/zaV0VcnvuuE1
yIge5DBM9vfqrc+vy3MV8Wd1bcVxSG97qf2BaucB7M+g15L99f/CAqNKLmTVBM/DfAw4XM3h4PPo
Ul48OcOmud+Yk74gDztEpjvHf2NqfmtVfjF82kDW13cHeEPz7RQekNCasAJH+LfbqAbGAAC8KnUM
1Jxoc8ddfLpjTbv9KtLfemUwQQ7eMx++qXoGn+wsej22jIPwPumvoTddftwtHbzR/N2I/4VjVCkm
PwUE9PkGM2g5KIwIo+ZUhtDzHrpsON6/4QL5zGPDOXVMnsbkNKsJ6oEWUyAMn6csu99M6HCYp7aw
LR9a0AP3Lpv3CEbcEXoEjcG/2UZWHL3t62w+ZrWe6rz/wKON3GgStPrK3Z92LLIQ7bJR8GkUA2Y4
FSHfeeQLyRLCQEZr431QHd0xtZunLoi/YxnROZxLSVl/WcWaMaZ9HRvlkE/yAM47IRBT32lNvX3N
Nt4W/Gsfz9tIM8F5Q2m0ysTqAOo+/yUgU9s9lOZ3DGoqRNOVPxri17Ar1bsf6uvVsZKsGpfelg3F
nidkpYrRJCpY5EIgS/Rbccid25s24YRSoTF68kHn1+RU/M3HejppJzJZLzPmM83RIgw3CUN3sUT8
WwQ8jfT0eZs9CwlBiS2NY8m6q2t7uknJ2QMvWds8vFA8+kCzbJgSnecze+r5grKIeY3BLqhiSAqA
L9CLq0Bp5EIDzUgkOfeUFs5iFE1jdVfR7plPXNb/8wngNsAaI8NxUna4rvW/lzjI8qHO3SOKrXfu
/kZTv5wllYRUfUqz9wBkSsPstdhydI6p146HOzjrmmoJ6PTfM4Fo/tacMLb3nl8FMsHtphzsw2Yc
Am1n6LMnkj3PxWKQZRtBH/rkUmlaUnR5ZpASLmGL47lccmQBX2/WgI582LuuJDjB2Ys02s/jMV+V
tSaNasTnBjrkYekcyhDf2OuSC/biIrOeB/ltbFFh+AyYkiOUSECoPitnvxK88bI1vPv3AkT4pjpA
D+F6X0DDN8h8Ol6jpWzZi3IlR8iSwgRffLa7Sm8tPcaR2na2ztUBnppVTPwxOQwJtgbV6PByzlXH
r2novPno7abQv7gprGphYw4jhLlxP7d+J6+2DCcqEchBhzLrGQ0qfRcaCCDtsF5HKDXy7U2MDVz4
HLQc5CwWbudtsjQUgzE3MwnXLB297fZzfAtVylFvaq9+6mbPKkm2VJqlohNf4JyU2D2+KgVAU3u+
oCJBZ5ew8dyPYnWqqeMhKRCq5DA0ffAx/1gCGj40Sn3TjFlzy5NvtCAE+N+L0CY9mWINLWXAiC6J
sttgye+paqwDokIIAmnw/ywFYz7zhF2lVG35JqEZX4fozMTbGE+nfk/dMntAvaER1Gm9x+Zif/Ze
3whJ46rdEc6Yg7PuxP9jkF04kxteD96YN286PfMV2OdpUR87UXqWLYnovUvLBPnm2xetpciM4Zcj
BO1uGMhK/4Y8Wzuw1tPimtc0ZUJDa43nkDw/mBgfh6/EqJ2sMGS5jWTITAOhkFsL3hkSvCo+hN0n
wYDgLUiEmVhoY7I8+oSb7XFWS+3pQiXisTop6+Bc0WWjrK6dKasdLrv9wsvQsapXontlffVqwALG
YeWhyEtOG6hyyOCs8KHbEwta4FEb4MhrxhLtj0HNNFPNVLCATS3A/KWy2dTUa5hGHDwgsj7PFUIr
9XZsaQgXY2DLnOSf6gFQJToIqmgM41Sqn/9gBpA9dPPS1UsERS1yRfSOM3OWJtxSnvGmYNWBteHP
asDXKMBtFEYMLCfWcR0bcZcANzxBNHot0Mx00Mtj1vplj5ZzCiKOW/zxRRXKr+R7tZ0fIPHxsCD/
4LBfGHXKHAACvH+v690caXiVCcRseKWmIOsgPGymq5MC91z7/SuMo1TVFpBIwFywbAwmpkfER6z+
S+ZhA9msYNTk098X+mmQyElV/iLcti9Z2ITPHWBl+5f9sWyCwn2uEYGupL+06Y9yTrwDBl8hecxz
XuStS9/pgHx4GmMYcyje2v3jBTjwADOuiLrGrQp5DHpsLV+Uh36obGTesy8ZCOcUOcbKuXn8uvIQ
3GyQxQF69EpmxYjxTNoGDmBssdUY3Kk8Xo0tlQTUdMBIhtG+nTuu59h/HT9O/eXmHuMakHxup9vb
3B69PfpoVkBwIeRWt0TCHcquzcY3NnCyeZz9Gcre/G8bWSs1G/NzLfHEajsu/V7C3YE2SHmXhfeg
htN5WtAaDpnX3mdAlYgd5StfblGsBBfm2sx/7x+ovqEk9DczX3rjeVNMi87HSIzlmlV4xyUTzUoc
QAzFvX/DbTocaINwSEDOq8UTlr1KiexG6ChYPzqZvESqteXUxegHiCND5zvXTTt3RY6l2XInKtjf
MyoQ8RpD6Rrkmeq9np1DlPe2bSXLfZ0FFbqUXN5e05IX38CkMdXZ0NiJTrbqKFS8u2sI5yg4sGRi
+lRHyxwOTGxqbmOL//Kciniqr/eMTL5kkMevHUqUnvqSiiPYJWI4di7aK7U1sh6Cc+7aFvCFt8QV
QIAkcBtSchnUVyfY5gzz/FsAtlV33MjwJ5fAYUNahip+IGAiRuMSTAKTXUQr/SU4gBNhE9FupaJC
yUEGQJsqaia2vBs2yZ9Gwv1fwXqkwy437WxA9q+EWoHV14bo6M5D2Rd64YPV9Unu7Ai5X6f3fGZr
EkRfA5vZeH2tqzJXt7nXOmWJcKi137KfxdexMDRi5/5qfT6RXuK70Zm6xHyLktRBSQrrMrEm1Xwr
AMfWZ1vhgXJrdrr1arYZ/4roGRYRkIIEqOV5ttazhBm20ubm+VVk2wogdBjRVN2aEQiz2AB9wTDm
Kdm/vGR8JgNTLHPri5ll2DdFjOVkBtuLIXonQTwtORtn73md2b4xMNI2hw5j79dTjVYILsX+fcxY
v63XciUAArB0D8bo+dHaT+tof140b0OTpW36cf61CAwTWfkw+s7D4u4WfjwLzXdeSkwLF2XJuG2y
OIfoXkVDLP1WM8Qettn5GCXvAFaTZJL4seVN79xzNje4PBbySFRfGBp7RMTm/3QuG4Wug+qAyZCJ
6mnBaJn4QYcq56BLpUtpNtHT9Jr58Cht7OvRf6EYCIrPkp/7fnMmTuyLWKIwj73D8ds9SIV/3BU1
d+ySMuG23objCXMGReIdkVPc1Tc3CdxzlMBl1UV3oZudql0QUpsBLjBcnIukZxCmeP1fyWTzuIKG
pU+d8Wu29DsrP9GxN7MZmPgpyx4Lbswxdh2//LwcL3+ofxqRveACoNFJ+LWASi05M0BCCgOS0mci
iZc5ixVuUAAnQri5wy6lDFh+4Hrwznkw2d57DQYHYAQ4CL8+AW1YscTMl8LZqBGdcFsOvA1DHq2a
2SHQ4hStq6+FdebUChEvSaUyQLScB6YlU5mfIB6V6bR42cx+RSrNZ4HiW2pNxM3o21e9EpvyqEFi
UH5NKmevXQyEt5yLRAAK0DeCoiKgRbiL6nAZ7z64dQJeul0HPdPdBCaFl0WtgTR8MD/kIUl31nQf
2kc8kSmTiGo89tqxJmeBiY6qZBU1jrSXbdB/+upwhAjumhWVSOQpyMjq6kJltMq1mRzNn3EmJYqA
8hSoxBhaePJhQF/M/Fpt8wlMQPrThBElCUqIHNOlOdI3PeMK5AVxNoaYZc8hco7Z/EiwfXzskvFA
NEu5v/ArD9OaWX7cZai7ywLU+1MUv4vYkmiXW2Hunv0HJexisBKaVMAUz1RKg5D417FxAORPfFZB
sRowVL5pL9m2madQ0btLDip3GxttjNJ0b/uXXyfixiVRDbCU9g8zZbUzFxfR9OdgH2by3qT80esq
CQs8c72ToXG5PjO+rcq/NT/VWrgSLUszvDsvyg3DgyK+uxoH6kzYRhclxDaiqEhl4BGgkTU5Uhzn
1sqZ5ayjjP8RIfswy3gr9ZBtlc0MTeqrNnpd0R5loQJW+NSnI4MQlQ/KNFivKz6tHQA62nI0djEj
WstbFfNca3Aj3VKZq3qdyVGvSib51LVZRMtXXUHhhUx5ekdyiSIswYsoKiV9sgLgrhTTDs7HnB92
FqzE2bQhByFNuxCWI4Ead7G4y1Wyq0QoG6QB96OOJhaIXwn6p/wxDEXBaSuONIcc5xTQ/N1+6Htm
uYl7uw4xMWrkXxWDOGswEhyKaH6gWItCv+IPBwJXd1icPPB6gOzSKOPhqZKPD7plQK8sszshDqkg
ofBuJmGFmDRJucVMVRXh85xyEfTroyOlf6MGUm/DXBY1rTevouK+HjmF9irJFh1vqiOCAmguKhBA
0bmjZ0fN97zjpT41oGC4yDhTkCTSoSs7rEIv/mTM5bhCK9S51UVyCA8Q+02WfojR1PItr03GXMlo
Mw0j7BRsUNUvUDUrPLqvw864Pltmy92grnoOiGM7J3hwKHVA6aa4gvECoYc4FGye094H8cQ2Yo0B
VZbOKYwn1fWnBYbIyjJJvGxeUK34PyuPyQ54PkhzTKUpwfTnXrfp3lPmsw/q4Ix8F+w7q+Jfe1dW
6JkTgJkUo5hVt369n3Cmq5946pNvKdaXhMvzyHDFcbAGgHqtOpZjmuws1oCIUo5aoNZClNixvX/M
Yat8lES/AdoLcYw4rTxZPlBW5ceQnkR8Hl4avD50YTfWRUCxkRaD1Lb7nwoG8Nj46xNbYyH+unyO
J7WfeWPdDpArc+LUPtc+rb/HOGGAJx49G48+TOzlBGy3iSn1eeBWlPCpgWkkXIxByjBDoyhNsW9c
GdHixcD0Jyba7oSdyQppmlk6Eo9i+uCwXoFo9q03v5H90/S9lXCU3NHE8SCyBghB4JiQqZwSv5Ku
BimVfDGkD/200KjprlDXenPr1mANJgKCQVPklGIDmWj066ySVHYUtsHAW2EauCUXhBnVb71Uy5qO
ij2+l50j+iGtZd/INqEvs+Npj18sDhjLDRnlk7W5398JsONkygWGyfcPY163g1rBnmvAusXAV2p8
VnHsndiKngZk9pEbcn1jRlW9rg4Tnr0NT/QsiXDy7BkAJjCl+BY4ZdwvxhifM8jGhk23wrlZqTMZ
RyElUufJDO0NyuSYFnxmpyMFT2U8hHVch2wPQnv2QE5yo0Q925UI2IPgpXmgKpWI/qwsVU0/nb1c
DgI6ixd8Puxk5s7BZkZ9mZ4pEIJCswrYyWtVu44GGuky875vOL6NQ0Bh0g903eI1E9g40M8rimG2
7idCSjI71ijMmZ0SAxkkl2ck+BglNlE9ijpcyd978sehAnOAPm6VG26TTITzah2GUD/fNhf15BHV
Upee31u2g90SQ0eNpVGSURwT6YoQycZdhwBmj3w8pVO6W3yUcNrrbguT2jFa5KyWuFqAT66udRrz
QFvGUYT6FMo/Ibgsrm/51QMUbGUYoaDoZPViZqc5sII7C6g/zbvRNyjiBPTBn4D0AarcSiljATBS
t4//UPiH+K+eAOr2yjP5yQNEtpNYj7u1I9M/bgG4RtYotdlkwGKxOv4dAZMBG1890wG1HgWGNWHF
79+iJA+1LWP1sFp3dccVrRxSy4IVhKDrhADWl11+TgEw7wWWCA91/GyzD7w6kkjOlv/5dvgTOLVp
ke72TmTmgmXa6SxwzXsAWcHaw4FeYn3T1MRpXbEBDnxr6D6Bf3go0SMgI/X2AgKd4BbeY2vtVzbF
ceROvpLl9x4MFBSIcmA/JKj5Urv6SYnKqtpk/kr29x1nIZGMi3+seGrP8TxqTmBYOn84hARLreGS
3AqiaCM9+i+TOwaHFJBiP2hgLYT51zkkF8+ZuvNcCZyHUGQY8KgN9Qvk/2fQoROgK+xRnUJN9LGT
jxwW2urMcGeGi5HVnonickIAOL8QZjmuokYSUxt2gLU2SzA70dA3xZJ2+HDml4kx863eBCMNTbs7
wyS5nqhgCLA226ybE6umMOMYg9Xg78VDRWPRHXjRS0H12tE54udB1ltjSTGdofSHRBxdR5GwEWJ5
EsZjSNRa35Y9D7yHZB0kt3D+VhiRveMJzqdnT8kPW0CZJ0LSM84tpOqqxTlTLuBdmlFmciLgUoeR
iS7fgPqvmWLjrKTOZhiOt8aBN89CCpL1FJlEkzASnHoR8oNZSKUzL0vwZCEke53A+jZkjVg2IqAp
Jt8zN3aIt0rW2Qe2Yv7Z93KI6LOhnmV3YyisUUNgo7Dc9J2Bj+ea6DjMW/fmn/BFjQGnEF02wwLC
+CPi0XBPw1SlQ9q1gUG1SYEjDyTMJZItBgq6//4mB5T7GqxR9V8aI3lxBM9Xzt8pAGJOjllB3DYH
CNo8g7t46zJowqwc0ovJ0D58ejZDW8wnIBd3Fe2bLlohFwgRg1WSikM8p4jvJyV2jJGpgAKJB84B
viD2SviCN9tB44t+BPwkHLL/JiL74YWW1UbXQzUPp/PY9u52i1Fqlshbw5FweCaujALiRa2XJOu5
z7h2/3WijlAXjIi673wIAK5zSXDqw5NH0caYH7KlrN7zONPqvldwbw9+N0+2NcTogIK+4VnPNW2z
DJ0vYMBeAIbu5VS+2yq5OPZP9xwtXtkzorFnEfLUKR154e3ajpgpWyJDeOashg39m1QMlhblGthx
I1EhGxi5TRLOtTphHK09ZWnD20QbPvXN2KTDqt1/F7Fl5Gqc783p/HGUruUc7KGcn2yJ1ofqcZ4h
Rz7LkGdGjBOiCXfrlHiV3Xj1ftRz/Tj2h5aDkPx1X66V+7o8jIFIhutypfrACArX09RGF01Erphc
3fjgJa/qMeHjkuX+Ck1zXXxAMg4JED0L5AOKjN//3BQk4gO2ymbWvXDgqjRcC4Ft7JB0evQLKvMk
enNSgFql4gBhKgjdMq1X3S4FljW/aiDG0zYzsIIFuCuaK/9OvT5ERW1KWbKu18IXFAAVAr7cB56m
uKBS1R8aFfS+0QaXcueNuMLmt37p6mdabk6aFQWbYZsnQs7JUBF5sEB+rpSgeUwWq8ixGWpa1ScA
8y6FoVSdgZx2oOCiC/TCfGGG5oZUTBfkquW5boW8GCqoT/MNa/3IDBVRs4yiJjrInqrSPGZ65z34
pLviiZZuBly+AJZqOEhuGYaHutBvTZHnPO1PAFY5zlMLRhMcUarFWhPZSoRElh9Bx7wf/Q8NPH0h
PlP5vsx0lKs7iY4rS+n6Wn+flQaBWFGjbb5r/VDWr4XiDP/pdxpvhDbhYIYez5lwuRtPfAo9rxLn
LKFREQ3DBi4ROkZlKQN3RqmKiL8Wg40QVQf0ilWF2NKyXkC7xkx2hPPFFTauynwt6DBgxjCt5YF5
/aXbN58WDMpDtsquLe2lTsoo4WuLB3yq/4OSCfI4j/y5r3tJkv3MPu96uEXJcdaUVls/cv0KwcYw
dz5C/6ml09OSKHWBbDDf9UJBAFlO+pq+thtw0LbA6LkznuR3bkDDeWxISo4ceThAHCfEokzvGLNz
na2GuFPKK84hUFOVi4I05lX7wAhD/HKrdtsiZxROydJtx7ozH/oGP5LshN6Zz6uSgYOYJQ9/OCxf
fp25YhvG4Y910iPc97Jy4YYyRHQoWcz4Pz4TKYgB4NTtz9HOzSKaPKPWEpwnvmYGmaHDtqxP8X7F
zcwKMaCq5crFjgf4WqRybwiHFuPTlRD5ZQ/CFjqAIHhGeCQ7MQfADkUuT9iR5OUO2MiH3f/ul/YK
d/97GWAoVnvdXHMU/K0u9ozw9wS/F63Iq0K4GsQZnh08A4OX6iQzjs73BSi6UwX/oE4I9PMzuSdT
zs9UNHB1ewVMSK2SspA8UfODzHzA/Nv0jVWIpIA33HyHackrutpOMF4cCRuS+O0cXxgY9caaTv8W
Bkf15woQz/keEndpENCDvhU2+wIhirVuXdFkgqb1Fz59mFRsSmp2mi5SKauwUKrd0gDkrgD5lN8B
aVpgxv/GRqAW66sV1ksP6nOOzJBgp9lJ96yq+1BrTEEuLICXCkGBZ7g9wT848FnJirYEleuOZ9U0
LTgyTEj4CdcrIYMcmj/+762wFwnCY8E7fSXWRMpMtkWCnaHpmXwnB9QZieyBP9gXcRUoo2eIiwj3
PJBCxJ+YI7BDlgo221W3IrkKwoY9WCzOeBPooWIKQ1Tquvs90hKCAmrWJZt27eYfd0esQI7QuQp/
XHK7PlM1Cvy1ltsL9jil26nwqz7T8KFXEXQmH6zf6IGUTXBznTvRoMbpGKVXdg/ieoo/uGPl9x+L
8vOSN1WmVH9xfpA+LjyTaNMgwW4y38MAsZE16tmwqRm6joMgtYsA3KAhI77vDCT2eBysGugnGjNO
azhOxTG6KjUj2MRcn8LYAOSCxbYNc6NmRw0ccr2XxDvZ+ap7aT4ugcHItBSRwZC5wTNtUAycPZwX
CRtz77G9ncTA38RdvfASSjtdV8C1TzRvb5jYg0lDZZLW4gV0X76pqjSx83eWjqCs8Qd/K4Zf2EpQ
r7hGI0TIRlpvtXwvTcWXiDl/x3XE6udHNtb4Vv0bmPNTQO1UZZUZjmlukYOiCsBDNBoyBdDWZZK/
6tmVpuub5rKR1FzsjVRI9N+RMS1Pr93EE//JeNF6eWcLD5jd96i6Noqop+ptPpR3rqf/zqsf2WL+
7qyowiVi+A5wD3xICGplU0chGC+8md9dd8xRNfIKugbYUi0OOHm6MgKkfbsSgGMdCInGyPM4zTf9
1JfFbUR5NUCfddkXZywN/PgtjidOD9tIuStozbMXtGBedQmHDAHaiQLgqPsX/xOrudLbExFL2Dvf
EU7dZ+0S8VsTzh1EaHc0EkeTqXWNL87j2Uz8zicJ3Bc0L0GYvbSk5TCQ/ji16t5d+zKjb5ycbK2/
bk0XFEL/TfVXOkkO1x/+Qagk8YxUz5rNvNZB3bbqLf33YyVXLT86jp3akuHwwU7Jwza6IcDJRu5V
WIH5+IF5PIF/sgBt1V/bJL2VGK+2nf/PHbgDBxEt9XTX4UVMu2sw9mwLIPHPNh9mbxAX69cfotFa
EZeoqGNyZcjQCDZuaovZzjBGSTD8ydrpUUJsXyMFJglx1t5vEYGuy5LYSNgV2NUyFCixRi06mJB7
rK2FvYpI/bWLSC9E4lyjEC9na45U5PuTopgkEkYAd1hU0zh0wydjkVPsigmPIpDS6GLFW/7RQ0Pn
vw3RSZ8L6sAYXguCZ0nTEC6dDAwxr18oVH0rwUL6Lnk+CmGCQyusnojPOrpDVmJ1mq3Z+DQbyx7U
3CwvQQ3zAkSa1hnOtY18r1bb+am0Ik8nbrbSK3aarbDImVmLF3nOdjG2VuXY4WAITnTmai3DzzYZ
6KWLtcgOccT2uKtrGjZpy3hhzR425Vj3ZVxtDOfbWM3+BCliZuBI0QrShjgpQSMG1eBQqIYumWc5
KGasHt/qT1jyYmwYC1saOOllheJVPVqs+ZNQzEYNqiBrQ3AKWVGlD0P3xt129zNieinx29NGF9X7
J6azpLNV1tpVoS3VAGnwGAdOq0Eo0f2Oq/iazYWxu2Hw75kpoCGfNas55KNCa/2Tyfgd6OVUA6aD
uxIdEUpJ20h8oNRyQPasOCAHsqKFtHNCuThAA1Zkr+WG9mAYq45bqZcMTz/ivcl1j/FGKPyHhDLU
qS/cN9LNLpm8tvR1JH2sHu1PbisaQKwFDuOfvaBefH9Tldk3XSpvpmPtArH2d0Eve+bI/Fc6Ui3i
ARAs3fkG/3xgBlQL9q2F4BJpEv9QgiX9PYKKOgzUw1O2KHMZkGt4RCUSfMpvWBA0pjYhEQUIokeM
pIEM+F9Z+c0fFAAKv8DJ3Igmxj7PPZLAKK5/8fYngwdOIt1gosZDiDtMRPr5QvIVul2bctUBlHUs
JHBLMckz4quO7GCGHM7FtPQcgtlmuPW0Mki/J2Tw1ukLE5y3v6jACitgQ6A9cSg2+78gQssA+qIo
ypag6doJuXKKg1pKsDHDfswLkW9+x5LpXmKPh29Ohk4s4rf71hI6Z315Ckfy7jYxJHOijJ4el/NP
OfEpQw0d+4Ujx1jyUJyyNmBhbNZf9Bvdb/l3AW/WT2RGjR5B/jXgR7PpEflrtDujxbdMIGghHvkt
/sAYTAGxTzWZY92rTouJ4qsXmtc9vFj7NIuk4s8zATbzkSOZLyaE6ljBUUmCm7pGEnUWcHTlb2cI
nm8xV4bI4wH3D+BwNPIFxT9IGrUW5snO7P78qzbUFT19SelVX8ZnKwf2imiWtyKw3fLEMhmpaAHb
3ePfwGoUC959XSxzAkn78gYZ+iCkP9keOfW0Q4OUQ3gQTkFdSEIl6gWa0nfFk4IaQBoonmKj7OrZ
a1Ug8nkQgVowMewg2+RK55wbv/eYxEJwy1alUvTyKhjl6aVisXklAxPJGr+s8fI7L/PCrDjlLtq3
cRWLJPBD3r/WLHaipv8JMmM54REs8aJMxCwXLlHnMzLAyAPY9qQNSgTDYrZajiEF4WUFOGNKMf5z
jDbBbU8kgdhWs9xI2O5nrkaRV6J3w7mBp2j3msZ6bF0gednXcqcGpj5BjgiIJr7KMXmdN5m9PbU/
ZLwdcoefeL9Ql2u7obdo+dRhxdVwN/dTZZsrcNmUg25vox/Jq0Wy5TC03IJdvWYglbHAcg47KVBz
nUatAq2PiqZhQ9n+dr7ShUMqmJMed+vQPj5rOCgtjh573gECsOYg/WPI4L0hiwt5Wuovno/lGxpp
gy5dXDa14fek13OhK00n1WcQRfB7SdETSIkb6mRjcKcFMs88IwyX8Ml9w6y/tQkJseCZr2Vgj7uB
wdaaJZtwkfneNUUO/RA1VLPMyQ7RfG73dJAXs9yz27/kfhEOSgmK7b1HPAgHRRbVnDDSMma7P6TI
OmX1VZVjK46T+LyWtT1ixES0juf4PyFuff25jbmY2GKlEebv0BBZNPHD/dj9BchE5yI/FP2rkKBz
QjoiJNs+ay1mYq+PRtqQTjIoMhsvHPV+2G4BKjcALl7oUR0phrXoMcgQNzXB32/OD5Vodkv76n30
uOsipaC3AIlT/vQvLp7iHaNcCdyeVlXRghVfpqwV6tLQuqz2KtDed5uK967TqL1locSfShJ7IfBZ
xaJmQtLG+XOcs2M82GlSFwcaEN+5dLVK5W8a3iRh2EE364XuhjtpvnfS5Kya/TgM3Jd+rDIjRfkI
inzmT4PUqHF/T4Ite2luEymD2EswiEGDTgB7Dz7vSHIQdXi6uKAthyifm4h0Nb196+xWWWX8KKLo
fUK5V+qgaP/lF66CT2HPQt9gWDsJ+AUnp7Jbg+9AGQCynhLPlCgh5n1rXb6ACcBk+96/I90EjU3X
4KVMufmZoxBtYQWSi3xGqtwEflrAB6BI5Xair+RoCYYz6aTFuHwl+NjsbAyi71btowHrianBZFJc
y5qf4P9BVUx3sIQiGrbHc+IewHKOpTKidzY3wBHokeAHtnDkDenPPprg2ArCpEZDsZcYT9wuPm9J
F7PJ7gmCSMODlWAk4+m1OK91FyJ39Yk62jFF/7vTZ6vVZe0kkZEd+2+QaBkya/mrB00xzOi2ZRgd
S7q8Lp9Rt1usL+D2UdMMOH0Px6REd9o/jIX001vnNHVCxCsDS3TnqLbHcDg355GMgrB6awDgIP+n
fsUzVrl9Z1gimxAE1bjqv4c1F7JNF6mi5EvwbKkugXofdiPMzijr1ichYTWT6h+Jkhy1rfnYKNws
wW6ZkdJSiludaRuoSOfAjtzh1zqRqfJAlARC5f4hK3L/QXDPYAyeuluO04yA2tTiUxXcwgOH3CeG
7NWU/Sv+wbW9gJaX2N9aTycx/cRg5xHDbhFus9SMEHWtoyD5SHLu0DwUEQiTHozJdXlKls8Ps4II
cHmRrSt2tnwmlNmZbGB1q5wNoEtNm6qU+7NfM4MJFD+uhWnnyZXP5bK7srBXboZmx7xNLNOPY/gN
Esy1hV3GSrK2AVwHHu0kOnYkUUFmmLIPNdJCMDO5LOE/OFzAMpCmh+aIQ9Byriu8qk2T0hzMe8db
Q6wU2JEnuZ1PjVL0rAU8Vmvjh/iXAbxiascc9mm3vzaq9hDQTZ/hEdujmbJ3exBopz0UY19KJQ3s
WMbJ5y1LyRiZ6K5ItKx8yiJh8meH9jgbawdz5h4vZb0BODTvgzBzqju/R45nBuLsXVbIFCnLTT83
x0dzL9mtHBVGlwbrqAPLZp/2lGW6tRDZCzWQjTYL9Vuwl8gibNDL/VBtmajIegr1d+R68GuT/I5h
ezHEo0BGPIeqt0y/OkaAkQ5V2T/QQ0FLwCctel3e7Fz6sHf0GHPltvwoTXGQ7l572ceAVUu2rUKT
aFniLtaC/G6jlO9/SC6hwMMZd3AdzHH+s4hhwjOpKVYEdt1ztQI15sI1L7ggBvtdLqYydrmodxFP
P8c0iRBx3yJjDNoQW95hs/R90F7QjJv+ZHcq2Itcp0baygjjfDJ9BynbatKYniW+MEHs2Xa30o7y
QEfI3A93ak+d3HD5X0dZ9HBxhdj/vcSpFUuiknLHc4Ov8esdq3uys2iV1czGRkJaAfTFhpHWG4Va
R0YloY6LrJ/Eh3Lnm79IZLgIEk63Tua+a1k5lGGczGJRP50fgnS37/+fKkZOERP8CEtREo0xG+f+
y3OIQUPA3/M24mLYKkTNQjADom+ExcEvt6SnL2UP0yvQad2fC3oA7UTXBjH+k+GP8YAfj6txCpiY
zDiGwPwWGhoH8rg4AlLkVA/ClX4XSW0OeWsfIniAEFiPljYlVqg+WNUdaVPyuK/bxLAHpGQEiCmE
BbPr/rdyXDZgUnDTHj57ywELNevUZwXCrjU3l8tGOSUHOGcCmXDuO6KBXp3iBYI943UZzEbifcaX
teHLn3xO+cuGXouAfWk3x7wyjB/rQ0LvC1Btj5SmoTn2Hm80pgl1zhPY0efbI78IzAogP6jK9SIf
mucJ8jKObvoA692YkWaNn1BL7hohQMwZens/ghmxgmlH8AcmnK1Kjhx4VVa3pc3/ionaA9B3zTbG
Bnb/RNE8klY2DPPacUGwdVZr/JMymycWaQ6ca/DmRmEXwb3w3ZP6UbdwdWBx+xDurQT7yqWwqPpC
WZZIBIuwyer+qLslGejoyFeZqQYhReGnuQYg4zgTT3ZodbciWUxLGSnkyq3zaQAOgooa5fSH68yC
FYXYId+vTHdXTFRFsqLYGnehBoFFkITUnzIGRvQHov2Yb8sRLPmqvaBetlVSfSHANK6loSG0Zzl7
Zr0KmyzpvZYGFJ+ypnqPc3jvAmSDWtIVw1GRQ7qbNcvomKzzOQ3P31QcquLc34Pp1VQxfXMD+tME
bZoikikesFM7wBvCxtJo5UCyXfkY6uppJ8MZIpfW0zELMAk6aVSQhBQxV+n9ouLifHvP6XdFGHs1
cULuz/kuFGEaESaegdxeDSTZoqK5GZnYFjvSq6qmnypLE8dckttSruU65dvT3QR62Qk2zUuTf0ea
58KLg6hTvRfH6ZBXCDLKk3LUOX9dX/h/xHdWWPgOK/viXdqwvN1wmEk+WIZFycQM8C8Q47K4pzSD
UGxBFqoymcoKWGZrAcYeYsjPU75u588Gz8FqrdxPiyQh1Bgvaf+OGsXmZgvDAQvNojNDufcteOos
/UkpxHQ7U0+JHWGnFg0HMOSGGI67al19tqZS422QYPcMQGr4v2lCoTthGE+OrrEVnbuladomDPPQ
r8Wy5YIN6hU0RYEn3ppoPnhQcYvJj8DwA1E+944r4T4VZBXuFozkAWvSKOpFN8o6qesGLD5mVr2r
DY3x3a+Y8tGZ39d+ltibWOVOk8tgGmrlLgc/xOgsbGG/YgG7gjZ+3o730kHtuozJGt0BnW5O75DY
pUs6En16zCcnkVg6VcAJF1W41jWTEqRVzUFi7NDeLqmm/dKE3JNS7m1sUZoKkxR6IzwYyuKHAPBO
QoUdRIcB4dph8NO+e7zb6sn6y7/SCNJsy/oI8ZN6RySlT02TjMuG7t/anPk1aaRoHLCiHYCX//af
RXZMEaFlvtHGTpEHUkzdIhdqyGgBqRomRFpkm4gYv9OC7ackgpjmS+qVQYW8GCrPTnJxa4ToWKky
BngB9KzJiSCTVGSrSZ9gM6O8sMNoDO5/qXvNGNZSIx5eX/6ZDC3brRoMjA/+xea8KIQvYQxWv+y/
e9f6jamE9T+UYM/faimLks4MQ0ANLIj0daF4o1oYa4zcwAC82QrSVPTVPOj0THShvTKmlJlGeWrw
8KPxylbfHMMV4kOwbLDxzSfViUDdGQw0h0lPjljSmLPSjADfH4idPg3Y9ujEsIWVhPnHQ5mtGiVN
hO3aEZcslO5No+Tv9hVy4FwiDYL31lHZWNKYGIIj5jKt2T7Hd32ngbF/qb0a6Iej4+FL45NJUkLu
JC6sGqx/28k/loFqYEUCjR6cffQOa3Mhp5l0t3i/z1isoBzlx+bLdrle7HSBlE3lrNByOMBbWNyX
jEZEkYoQQZjiNEBtCJFenHUlhx53c76RIOO89t4KH3x7jrDEauhxQInkA8r1Pvh2a4V/qh1cJmas
p/AH34vKT69ZWaJkC3p/eUEElXERVIFnWJs3UGgCis4E4Cw1qSHIPd+wx5iXqsEY6IGe5lYztExS
U56ceAD51vUg/xRdeU4zJxbdKd4u/G4Dl18PmGnmHyoK4SjeMA4FvfoZBC4I5LYIKtgOrdcp56li
08qzr+LMwYkLG7qHCTcdTUBVKGwsEBdaoE1fDMPq411DIMbyLS0+bEsCrfjykSJgAoLyabNs3upO
XiUafwGddjeRTK8yn1Rqg1T4V6pPh1rBH3egxdWJ6DPUpzt3Xh/VQ/vtzJHlUfhhB961ULv695i8
RQl1dwehaJgS5yB7l88uTQmXdxn7rZczco9tI664Htk3i7m95Ynsnybwm81OhqHKpbyrc19MNfjT
gjy1nk06h/Q17IbYHrbTXTjdItVBG6vKvzI6hovjQDP4OxgOCDbtjSEdqskdXGM8Fa4koGp18d9k
+akbRjb+JbouBTIaoax3BY+dkr0h+0/owU7XQgRae2wjYlUhe7Favkekjq8KG09XrZPb5DweYQns
1cPcmgfpNpP2POOGarW+jGXC/LxHpCW5pKHF5nFzTF2BsNzFZBOiEA2EGceGkIbwPDAnQRHiHGIr
bAwnfvPz29cT4xPIB3kquPdv7DeJ6aQOWmjIPvRa7JtNgvIaKNyP1RegL8dwxeACFJR+M3HJTp6m
i6iqbOnLM0gVzNACcq/rHF5JmZ7UQVHRUJLKDwO509/NtotgBfzTxmpsJRxFRDTTh25M5SRCzfvz
SQmIDAITWG8nyn2Wnpr1p65/CzjUMq77ip4eCZp2JQcy7uP7hp4kkGe1uqnKpMwMb+f/ZzohtZam
+MiizHfK+8F+7pIPzapKmYks5f/qeopUXAO4XJwG+dyRWluq/I0h6esgi/8nNpmrV4YrklTeD2Rg
0/Ljj7etQMzkCxA9/VyjI4BAi6JbPl7Wrdq63ZWsQCqT/Jq5W9lPFmZM3hVARs8WoEr1WVet5kbC
2DOtPjSb5+JMYmmb3/n9KIzBDWwuBkXKjuLjXwLFXUEXgvzdJcucQXFewpKolYZw0Ap/jTBHe+6W
Dw3/ZdudVQq7nAjjoZf3wOzK/BNKW6vBgN1A/jr/92n9thoz8OzN37bod77gY2gzSX2rTt8IG1I3
+Fvdt/PndS1UzbePeRS98Sqc744J0nYb563wJlpU1iQzjFCkdPNsLfifcadPSUObHbqZtiOyO3KD
XkBGVSf9i0kNmLhKwfVBXJGEmqAk8ZflY2161XYRdfq9/ZD5SAa3g9ceufeN/E43meQ2Vjh2/XRD
hzwVo1s8MpGVcHgae3l/YcTSKnqnuSth/vEX2uANdy4Pz9i69jCGzWXG/2kYZlrB08xFNoqL0NCb
sZKut1l/bN9y9mIB8xChyFkuN39LtoKzd0JsAw45uyYyVLvRMkDHx+eHY1OxBROCyB0dLBo71uEL
8Fy9dbGDbhlZb4ItHgjRZyAlpqqu7QMSZlXICYoIHl0IEWcpDmdEMkvS+e6FDDeNmGFnSjFxRGb6
/8nJnEIdT7UxKhpkuwELFkVqxd2Xirb5JdA9K62bFsxK0TlPWwwznt7jSdrfFa60FsSeQJdx5jAo
6DUwySlFE/0POdLcCuIGVsJ/2rAzew4o1PmLxC69g94gi/PzdRFZO7dVPssFRgNcNhaNXwuchwhv
r4IyZSVBITevBsJLQlooPCwIJ5qYA1d38F08dqgdyVwAPtBD/37WxQVi9F50wHu1VTFo/Q+aris6
Ik7QrRgPQJ0muh1vx2NEwzdHaflByaVJNXgeQeb9pjat7Omq7ker3xbCDwVR21sLw+0TC4jech+u
xfbwFOV6jLEUs4faBixIDdboa6KcCIKeAunImQPO8od0o8BU1D9NXYVHR4e0pcLueodecqOwlg80
sZurpGDTeLllkW7MwxWQ4cxc8mDb74KEJ8p+3a+gGcH+l8mpbYhbPj6RDNBYLrVyu+K/5WMhyWSL
z3r/iQQ8oY1RFqeG8B9AOGLp5Yiok2lRwmdH6oMmX2B92B9vMnJphR7oDfOTApS7TEKlwfqQD1nf
vnPZ98Bv4OZU1V0URfqurCNEJuPHofUH3DlqPt7KNGeSJCjAvDYK/hv3s5UjilxhpcilJTADzkmn
zi93A/N9KhVlsZs4oFKmKxAE3KDwjWix/OPYsNh1Sq6O54CLfF3VG8JlzRIsjMe7t4QDx7m2KsGy
gD2SBpvNnte85ijTbE2qMAGVN3JxIaAkthb9WBW4Ca/DSfw5pIbL6b04nPPeVC+sA/jntJjhPWWs
nR4ZhgO28ljtqu2spUxC43zZMNo+I3LMr4kqid26y800IspT9j93LoX3sPGgQ1V6s7ZsJSogv1ua
n836ZcqymxINuEr/7N4pgjHwQpzmPNOElLjE0e0O2/ocrAusSVaTBseoO/o/44QEgHyVW9pymwlV
OdCIl8zKTBQ13fF562QahcIfx22tT+di04TJo+uxXpD4gu5iO3GgeCkfhmUQpb2UeXzFQ/a+3q2v
QeAW2gAIUWbVqeuUFSIc6Dqa4hZYIcDv7D5WqKeUajlgQ3Ux1/PGBuFZmymxmufBhRa9ufExCvuW
7RPAmQepJgZ2hp8JU3rsBE3jhOZk2m55+JTnySnv3bmxDROdHTiQKsoWbht7UAj/DSMEHITah9hu
+lYK+2ufkkUF3GFehlbD1emnp7X23l13qZq3+V4BoV9H+TIx9z032M3SnKYLx/pQCct0f6yEWX5u
Z/plxD+VL4RGZnH0lMjaQ9KORlI9Gsw/5D/+iHUpnKhwi3Ft08VomHtk71Qo/nWw4+RMWxQnrz++
vDDHhm3MYqgdlwYh5W3RIv26cc8N4o/YuQhmCKHgohVHUZwzMJn13FiL3U8CQAe0VcF+Xgoc4pHN
vE/N2AM8CQvRwph90tuIuoiFTvXVL1nRS4p3XjDqcRZ4xokMeLLbX9pLVVxuPWZxNh4TWAvGqgWT
7idcQUOrbpIumbCp9XI1LfleJqd8oyYOZkhJ9Hfsf2KBQGo7xku0e6UhUqJGqByuq0BoaHdH0v8X
AiQfau+i9qLM+muOBbpIYGGmwgmFKls/GIPcjUQlrwBebyKCdxAT719LRxBzJFI0g+SqnKXn+L+C
SMRpIAN2mG4R4bXmllaQVe/uR4zywAHDkxcv4Ly+kjnORBUEHO5Cl9n+6qSvYudRybXpMBMubMtT
UPqfCAb+kv+FJlIo6kwJSLCs0qNGZM0d+AWElzwi1kANXiJxB4kNy9viQlgM8jaFJhqJBvgYs8+E
iOk3oMyZ/Gyrv3FvC3CUvWPL9FeMc62JdfAH/5FjJhvSOQiB+vncfqou7dNOmaYRHrPyADAfklYZ
abnijE3ZmHFNJDMaDzeVZf9sYwmbnu/JkurtD8rN2/8qon2JbrTNRCBaZfF8e9bcRXQvR8nU18gL
qhm3gRxy6xHwU3UlC5J1i61Uv5IJrUk4BK+9I9A2CHRmq2CAIEjO5OJllp0i43eTYkU6lCXIZ+uk
3x29dstg24asE0fQlDaX7v3aoIM/7ah7AMMKO3Ms0FuAQM7EdHrVWEHp4Wyvlg1TLghaEVlDZilQ
j7QfPyJ82IAywbt/UFeituGvcqYX7bu7hER0/5BYrjs4w0vCvmh7kvC/ATyqPveul588OzlKHRME
zAMN5Cdv5EWLrK31VKI+/Z7c3zGGmp9KZ3o1mrf8eenah8DQ4nXoYHwP6H8WsERhQkf0+UhHW2Ca
9VwZSmgHrBpJ94IKelQadarOTdwNhuKN6n3nUp99r0mOSZDmHP/aN4rqSKczzn5WAo4iPd2lsUWh
p5qm4MbqPH1wAPlP+7Svlk59jaBgEbdHeMwjlueoI3h5UFmFFYswMNVA5p+aIZO3d5QOP0AgqH9h
LFLsVL+ZAEkE60Ars66vTDUv/ByuPje3J26fxzHmNGbVjSoIWTEX1oDdIp+oVF8zmbIcIaE7r+SX
1JGShEF5j1h5WkVRU2gxInhvyJzOcOyurWshs0IMdSg2msatLb3G9pUNWntEuTSJU7r+vP7/cC5k
pR68phF4r8/qSW8wuKttsc+9KDwYx8p3LteTQs1lOn/Y8oOb/9rWmRQKhhbzc8nmrW2nExwPmSm9
kBZ7QP8L4vbDZDujhhczlFiyDsK6kd5psSt39mqlqPLEVOB2YSzszZKfjTs8e0e/04xQwIEvKZJO
s8zjdr9MdtezOxJvnQNFe+54oFOe/08YpXQpZgnAThN9GuuyLBo9c6G7pytbrpJIgsTYBV4VdtwG
eT7BeZdGtlVLq7itykloRB3Sz3x0N/GA5wdNHhrKA1Sp8HQMdJNUxcJOi5E5YoqBMZ7PTsgR7C4p
ejESzHJ2IvuonBS5W9G1nbxYk6ZRdONLD6m6Q9uy9dhZDODy6Pv8ZqTNR2J9YoZTIqM1ktTPXcQ4
zovG+y757P4qiFBpgIYcNMFy0GrWn+QkWEsVF/9/UhSxTHhWp+bkTI2LV79BVaPmlV1aJP7DFB6C
kebz32PtiA8KflnkFIF6q5VHVqqSdS6f6DNBfhXsJY2Hmc62CBUmCkXOpEk7WabCFLa/KP4aq0/U
LYRf6dPBhUemDtJVSNu1ULAUCrsE9d1SxxXG8IpMC/Ic6j+iD0FPjJMLSlNaseOncDJILYFyLJ2T
e0IjNoGcNOToDykrW2+kQuwcNWfPAzt7ehZpcg8Nb4ov2KKZBOtOWAn3yOV08KkGj2bca5FEENfQ
0PnqP111VPKJgPimlV8w3mLs5BHHWc3M09xhO9e1Zz4e9OK+uM92ayYfpcSUEoUbOQfWMrrlCZJ1
tnPgyzly3VorL+ksJuCv9uhOPKXdQOuDVkn+iSl3nz/aawi/N5KyEz5U0FApLNOdK02rtAl5VIPS
W6F5lP0EZkqiuwReZ2wkZwaUUJxoVWYcx0KY0oScEt9HLEy+aZH634mALBzk3907KrwP9A/sj5qP
Me/5GjA6jRlQtbC2r1+4eQJ1hqnZJf9UwDYvrzWPT0u7WEV6Zw7ucHGVKc+KP8UoKZocvPMhkNid
QhKWGircB90micvyxQ3n0NWAA2GVfW/crbjEkossIcjW0Lqlav0I3UsrAymGcBCHTBVsu+YQgu3o
OUsIpULerhzaHUs+/P3EPd2k6AterDnYpRX/hpGNcKl3kIEfZ2gXeKqvFRKVM4JIn2USWXZM2UvO
pTghy3FVxUVCz8Y2OXHeeEkrAoig6tbnAWYXSDct5kG8Z5zpceFMD76UwzMBodKqULaFg4oWMgO9
x7hOKAw+qP8Dt5/IteIObeh0xvfYdSEHewctiIgk76REq+LqvGMs9wMceoBO31G1/J4P66frvv7o
GrfZrYJihfhxu5x2eKzjQLWIXBdMjRPiS1cgJ4Q/fJfy2nIjmTSYgtYSzCrfs4urEIqZfrtxCjxj
RJ9LZhSqCnz/oUn3P1uD6VlvICOn4qhx9I2bWoAPTdPvUy3kKLW99FkgY3X9YEZ8DhByJt5nnD6i
U9F6rB2Ky2g6fFcGzRwHlfWlvs3JRNh0o7B8JfA6141paLJbk7+CPgPyPedC5RIfP1sIKIishxce
mNoGYrlgZQMg0HORqozxiIe3ObtybOygTISV+M+kO3TygBqcIDTtkj3ZwzGSJBRd+p7PaVQAS7bl
ruB2h2oHyJZRyeuSd3GWSk8CqwDYtPzyLr1CVUDb5Kl/of6tc86zcPV9KzGfNVpjPzL+rbWCEhMb
VnY6bWmzW+VjSdTjt8fXR95rhnIiS5nYnrTkSdbOQNdmLH7aGSDg+SAkOCrORmI2dwDNMDMM1Lk0
zu1cXmh4IRlSd923qnRGBrUSDhBWAzSlBmXvGW4BCwHe5ZIj4qXsbQP2/MCyhDkWOmOWDLZeGiWT
r6UPfQg2jpSXID98yAiFYKfkI0xQMZyIoIqoJwTinuOcywnJqSea7TixIwYQgsNS1IW6FQBYxvo9
fHFby8FJUvYxZHFigY0BmF9FaCbJIJhFhv6v1XktI9JaLyiVI9lX4XjRPjDElQoEkIRs7tzFX5hP
2AD1aGlFCriSWXGP6zNo6/6XNPPQLwC+sCyzA95Ev/g6JMn/Z78ff59sbveev4ioAhGvVjofJhrj
mEfX7Xr5usJWWfWLiTDrzrrCG7QS951McpTgu+f6WzyFekbPjZkwdCK8VyRCILwxiZJQoW4DphHi
GgySzniS9RTt6oXko9tGceqwOy7INoFZIIbvYIVtLywrofcT5w0RBLa2vgZX3vhJ0Vb6DBzp7IjK
sferWrQspyqFQHy9iRVqlIIyinqBFeuOINRAL751Fw27CpTDwbPecWNDzrK3ip8NaUck5Y3OlPt8
mv3z9rWdegakYYfJGJ8ARlHEMhqFHOBmgkM/LrRPwf2WAWoqsRcmrO6CjJTSrSvELW/Ix/+5jNxF
Cj+Sv0SYiOjLwOthgsooxUJ8hZw36W65IyH9q6qWbtLhGILnFaQHG7MOaYRi0HAgj+wuwuRStqpo
Jo7R6m5VFbZyUwMsu+/LscY6uEcl9SUVAxbpflH6ACSvZE4W/SyXEY9ikXHWMhinJq58Oe/FtI/z
TJScOfk4Bd/GjWM0AQ1F60bFbs6Pna1a8M1HkHpTNTha6LMUbmIVRzNIGAI/3sAK3/65wa6izACk
iERlA83M2Tln6z6ib16q1g7Dsc6Jgwtk0w2kAph+9L3a//C7dg8DrSxVKa36fBWx8HH2YfyEv4eh
zL9QwJUJEV1FsPE3Bhd500sA5JhGXos7/7l9MOyWOfl3OsC7tAJc0kWWM7FIt1UB9zeIZYNjU19R
w1TTtQUEirKMsEk6AAuPwsqURHLThf3Q+Fun3E1dVHraZnHduvqfBJyh6tvzD65DCghieUV/uA6h
fZhZL1Y1yKc1CpgFUzlO3td+7WOW8vp4Ui+L8i1PDkKOC+Tg9CeAEQ0b9HUDVbKcNOpG972J6dOl
WDriupoHX1pwqh273gjdgj6+k0Y7MPNDVG/nsVp1sYAg7FG1tUWEdBk5XTLhgKwssdSxbKd3ubgN
bOMuGoysaG2s8U7agkcg7JFG8EKt2abPZXpz/HBToydbk1/FWs0/Ipt4t+h9XjYJf8dbcjbfXd6s
89nDQJkJYIs8DTVmW1p3P7LZIjVc2q5Rg2/xRAvbG9yLjaP4CCrh0Y/Mkk3cazhal3UVz8umCDMV
7G4SmeVz+D4FFYqzeaiqov67PNRIg0hbcHtKIyBtGC0furt+x/xiWfTIHLbGan3Z2dLX7mvD4p1S
/t6xLINvRO42Y5MKxK+pTWxL/rMKeVPD26/3p5JrNrIaxGMtTocIJwGVjFIFihAA5fyLRS0+5Ik9
yI8zl9TpVPNKC+iFbW/pmFdyVqGiFSIQzZKovIQ1H3QpvEAhCPvHIQM91H2eVB5ZMzs/QsqBqrno
Hq6ySgj6MJ48jazdCm3TkZMCmR/KZkNKWAK9YGsk44hegVKZShkif2iHEaA9/kHS8wOSeM6zpY1U
ExM9NBmODfDMxxmx3DI+EAaWu7AtFGDCgNGoxQcroYS9xkM+0U91IqXkU5CALTWvT2ARS3D9O5ev
pnfPmLdEKJntocJGZ5/qUWlmRWOLU19b1hfCxd5LXDLn0TyCrl7YmV7pXo2h/G3ykyiae0Mr+s6J
kbWdeiGSyAld4ifHxiDjSIPUTP8+gobTSVOZys3rC3vw7R+nRSqYiDgRp/4OuNRR4U3CsKJmxTVG
agJZBesspwP7FwwDlLx1r4uy6E5Vtrb0AWXfbUylLCorjjqVwCjVl+tChDGZg9QPeM0H5gTzCxOb
bK4r76V3Kw+FpLAgpcsUhHc5sT5ue269dhIWeFpg78CiSvnfvPUs99yKaKt2AZK5fUU0X05wV+tZ
ZeUsDzC/TLARBgTTI7oexJcnZvfyFDQZ9lgSk+P4We46w/ZfOE2kB1805/qtaB7R6msrSTl4eL+I
s+hbyFeqw2J7j7VKKsuTlokXmg2iZFit0JYHdX7mmPFYzTK7MROLcD4Z5Idb0VACngK8Ln3sjPXJ
v6bMqJ7dAwLEAIxGUQj9I0kApeHYoylDK2kFYSm0aJATTPb6L6yyeJh48B5s/VhydC0309ezY8p6
ZknjlMyshjjzInxIaFghn3Ttg4s3D2jd7RwChia9eraZcP5mStKWpJ7GaYYk7uKdtNDURdQYZ6ZT
2xxNtz27a7wZ9eToyIIXaGgpY7V1foSHy/M1I5qoxW2SD5EeyOpKam8Vz5oAsU1tlZ4kWOPW8Z8i
ebXN7LPVVUQt3/AS7cPbuNEx55NEoZeCKcZ4wlwgjfWCVm0tLiVio6VPTV0JtIAXmvdxphYJ8hEV
Y6jwTFiEzXjrb7FRrTLOCrCrEVG0UwJze8XUKZ4fzm5gSIKKM/xSrRwR4a1gZ5L4IUod1/KNJuQG
eurm0NOE6SZcF99ULfOnERFr8oHFhSJ48vqIt2puaKG5mKjR74n/kusowCpMbRwkHdh1XpBMHwl1
o7f2wFrKky8AfnZOFPX0yNIvtf0b+ZmBgX0p97r+aalir4Wqz7f1u5cGZuHX89UJDLAXcp5aeAfA
lNx2Lu2Cz3rZiANObdNsILVv+WtVOA81zf7z1hYGYlGiwwhxZFhZxVn5MBbDJcCPglu+4n0gUKIY
7pUOxUaPKGLIEbxwDDl4YNz5v+fDtome5EzXHL1wACHpNk/Hw1BqMamEpEDW5GjrvXDkF0dhHlr8
1pu6aeRMarQVPkvxviOpxt5kUC8mDT5SYjzwr6J7QjN50SSkajakTBxTz4cMzsMRl1fk38YqJX2d
TjCsVbEX9EYNCn6JTygMqAZBQ5FNGIifDOjfINaELXPu5tKxsni9a4Q2pIclItcFYPT4vyfKqMgO
izmSPJhOKP4nuTtm6yEHmNCsMH9m4fwiV0FNXlQdMYDWMVMdoUn4/SnEOHazFmXyYDnY89ML8V0D
7Z7Fxvud6bbt7VKDBf5BJmOuHAHrzzNNdL0Se16bvF/ePOqpp60sHt+jlUFeCYII5PF4l8WiCawe
XLh6lzSWYHnuoKmf6RbXVTiDtWxhm4ATruTfhHNhGvvssHvls8ds+91jwNyZ10E1kSEpIiXUoLDN
5fCQFjwM6m/SNYatOI3cTcvQalQYCsNEQiEgLOP9z0dcBRw+snTPgevWhTsOpc0NrJNSwXRGZDDi
7zAxmLXmDIUyU+OMvXGHi5XJpy49+G2O1nMatXRC1XMXpAjnE8Rs0Kb19jubhxrdlPQPlyffCO9V
Uc9v9xef8WOGjCE3FdMmfDUZVWcShzg/dSoTpROxKKejtZPy036LpK4687Om9piKvLINlxxkb2OP
7J26Q6Cv7+ElaPHnE8XZleIKA6xe2IIdAu+Fr1u62cSr5nOs3vLWY19BBtQxb2rzpyU4xir+aWxE
8orWksuXEsrgwD1lLZniLE/B2OMjy2NhMBMgEgOoP2LXt7dkLPhwwieBytsM/CVmUEDBQ0DLPAwv
f3auptXIQYax6Rh5xRtjN+UiMIo5V65yxPT0PBG1tjYAdVtLaR4C175Hlnqun+JvHFXZuOGobkrB
cnjccnNCPZ33Cq92OoqRHsd+Ev0b8+7EPXhAy4eakzMY9maq13GJPnKRshUVg0QF3CKqm5pCFhVa
+D7DKX3+WnYYltXkIGR98eCEVBphhNX5BEsReHBMew25bKqT+pgaGYGdwIK5iDpN0VF+rcrm84Yx
nXlYjWQbhAPm6uzLKJxGdfHvXlX9BYuowo5NndgKOD3A5Cs6ZyvwbQcNZiBo5c4oROixJ+6Aogb3
1VXh5RFhne2EiB21tplec70C7fnpkBXAYgj9QI2g8waKkiz5SgvDrBJ0U13TuQVIhLfDrjd8Pcp4
VCLiDOgtU3780RKK8cPFb2omLARW09A3mvqZRdljGHj3heKU1Rxc9zgg9ADII1tvMMvWkfcWi+7c
J/W0QjQ6QpIi1MvDv7w3eLgCXdUCLOHnYecbS0lxuEPv2TSUgFIqgDMsWjwSkAZT2jJgWs14o+2v
B/CTsbtpRyYR2uVLh+DBTazL6cbN2L8bWB0viqdPKPhpLfuJEGpNQXMvwypER6nA4xHhEa7Q2gCh
cGQb7I4yXrvTZm9UWF8rAT3GPxmPVp5HMpDF68hMjCoNnOo97Tle5au7SJM0HKe17hV6g0lLeLur
EgTD6CmqGTeAxEvGuoaU4bGykjewwY+haQMBu8nXHyeERHH51vyNt/RgIf8xaCMKyGudRX08RBHs
tVCQ63AxXSTAGN4ZW7kdvEfaa13+fVFj4BrE1nXP5cCsEJv9fjDy7s548i15NJ/nS6DzlfLprFIJ
vZfBeB4/XR2EBsVohzIWJsa1+xxLEdRgre9mCzvXB2K/A+xJEX33/1Y69W5fK3tB2u94kZw4AxMB
cnxwbZGEvy9Q7CwX3SoN9N+sk9xPHooO5xFooFmZgMmJh/tOzyEwIpyH/xX6dQfRZ1PCVvdUP3QB
hkKbAbOkUijeTnkKafhfoUkjIK1J6dRSVzXMuCcv+TxmbrkfAW/Q+qBVP2lGZKdLAmke77E6mFvT
xV+wfosNAOfQTAwIZTYBraLf39lEgUjnxSZGgaeDWNDLQemuX2CP+YKbi0LHI2swazwSUCYpm/K7
bf/fXboYVZ7IXruHcW8Qd3Nzoe6oiOPH0NXT7oGwgZS07OEtCfn+qDn3rPv6ems4q0F7xTHpgvWp
VgqY3u4900DGVBEb7U6NXRoSWKtfuiDY2P68AmAkYPLdPwCbUMHzKMd50SEPHk0TVk3YCOmMCrqp
/IBRfYQwBj4s9hsbqLJ0PdM57b7hhCF4HoH3k6czTag+cfRdPMBaRwVw+aCReuv6D29bgofFl2Q0
iYNaXWFCAXd52uTgVkAwV4yg/8e+pxckT7GgE/WjJh7p4uTdSovQJ3ASyAflBQr1fHmDLi4iaqL3
Mvg82uV9LrFS6a6vhRSKjSp+FUJ1KQqRIczq1zfLFwNNzE91KJNDwOJFM8N2PmX/KiF5bPS/lqnY
jr6JjPtZ0BdxqogrgGE3Pu+41ADyH7Za4ezhF7etnaXeU82Xe4WzJnBStE7erFweqew7XiYKZP2B
RY61hM0zT67xFY+aqVjB+FBIHdpI4n8247uKbl3zK8k9kWGay7Oy0n13TfoazkROBMaYIA1gPd29
DLawashY816TZM3NIgCzGWmfPk1k4UxovIYWVnL+N2RZfes3iGNJVKoJmyFpOKOaYjLzaME3LE7f
xNMB9ZCAKgPbT7Pcn6FVhpoGL7MarI8B/HuzrOUV1cye8VgzH+S7xYxs4iSKA+byme7l3LX8W6w+
E6h8w9aBi5A2Tv5su1Sifv/8AdD+BWmKsEGHO38SLSWjKNOlQXOWFZEXFLK28T8qbBjcgHmJ/WhP
Skqdb1d5RyublTC/nOCrGm6P5j1rYEwbqgJ3+OMpvbZieZEwVVTjJLF4gckOE/70nVZDYaR9Losu
v2VcaOHGFZcuoZkR95hR4k6puZMHza8sHathHg7y5UZzUPJepEI8IIahDnrYSoS5NPv2lHhGXyas
oJygnPyc0zmotlG8f/pxX5aKM5JwMut+afJdpL2sKEtg43EgkePAzs1uBzlHpi2zJ+8chtDRaoc7
ZtVn1DfNg4FGUBtFRrMerbKfowNW2FfBG9FbjhnTo7jeJXT+bjGqrb5/s69SWec8NZGLt8dJwwIt
CUPwR5ttYL6g8vBy9AL/Bcz9EuItQIiBI6ZURs1klFn5ScM8SGNahBOAYUvgETY0XxPQtBud1r1I
9eQowZMPb8rXMRDSItJ9LgOsYz2pzH1PQNdR9pLQSw+3BlcS693zF2qJJWrJGftQQpZIDdthdUw4
Ue8T8qLOjQuLSaYU2Dltaft2Prwt2ZruvfqCX2aCfcgN6CpCouw8sPAUzWS2EISdXabpxplSaChE
Gmx0vBlrFR6AcoP1hhScWtJbWTIH2ECmEG6e0OAcnLik1tvhxRHs7w3EsIIfPFLEYEZAXouzxls5
bwjPxHBG8hQVNWyw3nvk3aWBQkkwRA2G2J4p8phURymg5f49eJDrSA5SXZgGEuQBAsXiPKLGILyy
s8fcn0Mhy76ndO/QlBAkiChGFzfuitI/TZB8DFSbHUl5MgxRJeOl+Jn56CG5tXsUO+z2YWkIkCch
hRYGLtMSw3Lelh2KyoJ4Dqnn92qKPrDiphvFNU0vMNKYEKMdZyoND3NLm59ReKIK4X1Afa1fCooZ
B3eDdL9bGQdpmdG2NoI6YznfXKW/6C3I0at3GzOoUb5GLwOEiw1xhQBu8OlNujwIqazHzdDYBoEX
DnnxOIaJnCOFmrAKZ4XlmNfrW1z1WMuZ7K3KKtNMjz8w6hyLLKP0iZelougmW1yO4AVuwhLoKdsV
IBg/sETs9/PC+5hYGNLt5HHCkWxyKVVoA7lMLOlbG6x+OHBZV/NusAViUnwGs4Xcq+1DEru+X/eu
OfEoohfkc/4cPmTXFzcpPhn6AJ1O7NQMLxdSbbxmGNPSaWs37EppDC2XaUebLAXX8DDD1jSBQJ+o
NWe76WAUMZrRhRMpzIJJtq2DGiFcYZAxkPnSvHdzvDB3t186drDix4M3TrUydc7kXtvNT2iCJViu
7FAwsb9d6CsCxLFbQkWlpN3sZdLgardeoQbFdw+FNZOvfc7aFHaxLbAAYIS8+KIw7EgJSMpvNi8f
Mc6y8HNLD+pi/1tvB2R+/JMFYMntV13ctJC6nO5jrxmtM8YPp51jZ7JtfQ8KY4yn7pHd3lrtMMvu
kGU+fbALn/Le2MTP9ZH3cYXHJn6D1h3fy2k0H7xUsrM2HBH+Cm+kHta/HpSq1w4kzSdhU++69XSg
8yEcd9k2nS4h9G6SdNvpk5nFpBsJaSeOxEtWPqwyh/KUfPJnOV+3tDUiufQYH03CsqrJxjcpRRkc
vI4JlYvwwvGOE+Y6CCyfucwOrJSmNvNeETddg/TNVstbhK/VKdBA/4oXnZ7avng1yRHweHWzRiub
nMMYyUVtSiInO7U2Pj3lTB7+btBXhYaWbk/z28S98e6Ua8qhtvf+iYMgRTTr0YoUBbcZ/Yiz/y1W
LbOdcClNX5cw5wJ2Lv8WryKNJcqcukdCwPgLYNmgyml1bYQu4gNo+/GsZywiGHoatiYsE5/ixJar
KvdjdmgThlhqxpBaBkLmj94g8UmSopLAfjzHZFbPHl+IV7KKytknvFchP9erwu7IVoEuoEsbVuTG
5pl/MUeXmUnYbC8JYHHOO87WNYawHDrS6piuZUY2KGYuirO0rVy3Skbu6/NwJsBuJEc/4z6s+3Jg
OQFp0WhhU48Nq47pJjX+MM5OjOLz6/djO0Qh0cB4dNjLxMm3I5JedLtRj0YGAsnJmGOPnOKB3Zzd
LKf8v8DLiNqN8EzHq5LC4uAJODUh59rfA6PqWVnO7EKOZu8p9nNvDbILFUClaV0jj1ZRCMvRfcxE
ECzpLPFI+nqkNpNTD3al/9j2VhbnjT9tTvtkxtVQV5LF6BlPDfym2DYcua/HnD/IftsI11XSC91J
h6pdhNi82d2pM+qlJfGejnu9RVfsyx9090mmzfkORFEn/Vf1MQm4Zbkp7mVc3cJMIsIzDGoUisuB
kn+q2ioiACQwu0tUyADT8CAT/+1+xbrkZ9bhKPkFdUjvCMX53ULO3TdbKNEdXGw3OaLE9kt0d8/m
+UpXPBA2gbuJZa5AtdXJiHaTurZivIoZX4IMbe+Ue136soQdIVCDhc0upL6U4rOmdpYYuT7sHmSv
1v8Ocah85WL97agiAOVJAhxJs2bg4Grb3+z3HQSW/KqeqxxA1qlL1360OjQaD9HaImrVt4jfei7q
5PPGqLM/8cYlc3fawjEzOZRTsouHm8MbrXb6udxGyi7YjRcw/sZ4jAklT/XKqbTZLFSeQh5LCmRk
mhPZBO1jaW9qyEo78imdFaJEuhiKIqhrVSYKLJKu5oDjQ1dVIjkyDYN0jqadRf+POXBqQfQ7TkJG
F2dE+0OGLt5qMIHU94CszNV8WY7PiJi0FuQzrPGpgaA9BIOMFM8AUkjIhj0Xvl7KTvboXS2nFO4R
Zs0mg1Y4CVLnRprjmmXGGiAk9JoGYnaIwg0o/KJuw93Dx2GJMwqeko3z8Vs7AE3xqrlRd0Ih6VSx
1OXhefdAnK73QRHV/4H/4d5rcEtUa/qTAlkeRb83fG+mNUM70EF7RrxudU+2LKDPuxFGcPLvQdI4
D8YAo1TmbnHkgAfZa/LVx7Zj6ASzadMWMc9vkg9rATZJuTNdnFhEW1N+pajsEETDslxhbEJ1h4Ej
lZV6SqUk7/+htN6CXL+S7e4ax7jryXoSZsFdlISEi+yTrT0J4MbOoBSHWQx+aRDpYWgb7cvBgZ9A
Fk9wMsv64ZZHwT4rK/J27W/XRkbjY2Sxn6byTzrg4mDP1jp+BbBolZROEI3HLgyj3ybmrc+E1kH/
dlG3MFrXdauZ3rgF/oDX2gf4zWOcymQ3oK7Yvtssit5RVRvzEmwjs3lgulo3HVdvEc7NENocqNA+
Co7DkhaUNz0qc9pmvcPH6kmphhJKS8nRuc/jsOuASSVLzHiPFgSAiiFHIrQYkMZtFNmEVSB7/7mj
kRwOxDNgngkgIEFNwNnWV73+mlfr+P6TuorvYkqzMyBQkTNC/DEbpRCXLZgE+ZhQWOQE5pb87SoL
4XwSS4kRMYip/jvSYAZerCMvs2OZoSHGVOrJ8XGa7v+HIDplGngYQlv5duR9FpPgNUTG32F6dFzj
kKijDPgOIDclhQU5CqClYFRs87qKrSLSpAYY3KNB6i5CqwPdLUNz2/ZVMVsUm+dHy6z/lL/YKMw+
5GoFWRC5ayTM/rXkcium4rLCRdmZTelv1KRpoFAjDhDYTS44nYetqb9vcj/8l65bWxKOhEdgXVz6
CzvnMvsjkSOetT0KNxzekHY0wFdC9qiEvc+QEYCsu4iQj46XurzfivX6QjUlB2mBcTlsGYGSwosh
jMQmp9+nj4czTAAcDmm9JS+lYyQd5yJpUhlNhgiiibNoWNwUUhWwjwQIU9hB00JKUzB35GI7pNnE
uSdeOrKWzq32l8wr6ikJCZnNHw3xx3RW4IDRdE89hgri3LfNNRInO6m9zjr7P69agdv3/71U54nH
rncI5WWRNBjxQZz3NltAsI7/s0NK+H9diNcWQtKzIoYezZjCAtJl0JIexCn1TZ5hg4aFFA1bx8+X
N+mG2roKpSQaV+NNyh/QC3jBMjpT3dqS+4WqBRcXd6bBJM/yc8EyobM4/myTtHjPCYpT32fyWchE
j9BMUjriBRmX3AKcZ9G222OiiHiXwlxteP6Xmygo66y51XYMjDSRMcpZv1KkXQ4GaYcKxVkXLZPO
t78B5zayz0UfHthmnoT42XikUFhdAOFcmcNSiRdeWB6KcKdpgT2lXFjDxE3kr3O5Hc8h1XRF5Mkx
a81WnM5iq76OFL5LKfJ+tStHSLpI0Mqf2UWIfUOST9dNg7F50asN+VzbcwYwzNIV1X+zXJkNwlxG
RWiv0muWcVED4RHLbqifIlAHermUS2TodM7+QVFTkVkOqpo/UCnZfFBTHv6pCjmtywZQyj3dPBYL
JWFjga13vPHuMC+6/Vk/qS+IeuMxZ941RmU2MrjL7UO4fD2lafgYWxTSqNvYOffzMIFkqwBpKibm
0JUnEy6z4UMuzVsXAMZWN0CrJtIkBR/Kr7zYgStCA3+u7hWKcUXhXVKtUU2LMMRJujHHTz2P2CFY
o68ZBtiPWL5FMUF+cTo3/t7Be4DhD6CjZRYS2sgCeMwHuJyPx8fN43sYoxnXItfowyDJYoP9WRq2
TJad7uzKIDixYM/e+MzaSGQNWtcnZbSoWvi3N4vlaqoMSCIhtsJwT/rSn2xVreWe0yFXfCaOxfcr
oIko6jo1/3Fd9S5mWiO8Wl7bmQIZVKTHmh5L/PIUaJYRMS/C3mR2dOy/6pVLkpcU1+0wOx0p9eQt
HC33NxzGRg5SGVBwUjO7djAZssCNj3+rp0Fgrm1BxyRt+ulcv5JO45id23NCiNltbmWdOe887dqI
59ZrKmI2IIkS758AACIq0nZcV2MYs1Fm7MriNDmeexVLF6piTs/KDepgnYmP2Tg2EMOcqGzWnJMW
GyTFYKdKlScymgCRLcJJRKUNjfgwlXr6gHa54F3MHYBi6YA0QMtOfxU8IExSsbIQ1m46LjlZQY6E
IqUWJAPQ/jxYAlIe0vWRu9//MxZao7r9Q0ezYLUEYnu8LAOgjxUA1yINFT72vZmIGszZ/QxgK38f
DywiMoU0aWxOchlndJN+3mXDDbJrfwo6IzpPwIuUCIxmgZ7CWslrrN80X9Itl/aFUW08SOhpziro
pykHvQVoLMtwsWMVZf66cwWHb7Ydo9d6wOETGXFc8E46efa+gZ1qmR8hLWLVBNP3/ZqN/cEe924M
yeGIWvb9sYlbQ85IKRuW95/C3+ZqoFgTau5ntQwynueuXplINfhzKhMEXzcMBW9SYCSR9cGvCpIp
Lq4tjVDR38eqq+h4+jPIg/soN7JKwfDYnesehLB7BzVdMrve7yEIdB90c+P12K/lvxS02/yyHUX1
0BRWzNtR5cQFA4M++sxlejDPLfQdD5rd0Cc+7190/KH1LzuZiBEZPHJ9JNMXmfgcOEkgQ37+HQOS
oEw6zjoi9UJtVkJyBxuHWHCuybvye9/cq6nu6HMjaY3FDJTgk+yYZCDRdpEgzDBBMPwoQguhcAox
Hnixa2kroP7D5s4ZSw0DP0Bt7l//JZTaIMBXkgstTDEoXQIi6tS7hIHyQsWOXHLmnchB15sFPNle
qR9cn6VUIRPTJjpj2zZtS+EJSBbE0sxIkUFpHb+vhdKpNOWyLRPvJFkoHv7tDFB2yg4aFQSzsD2Q
E4bFKxFA3JvBozQBmx7qzO1Xrun6IiybGrYRA0Fk45eRPrw3Zk0tGpjIfNVjRVSlH9aYJruct4zd
6cGQxE/Anu2nyfGCVeuoNqpHrZ7of47ro9aqATr4EcRFyUM9fW1zmV7ZEcykyh69NM0zZZ58N2YN
hMZ3Z2zZcWg8IfYC5A9PYPndRWM5lbUkmZTEQMyfbTipyZEK6iJFS3v1kOG/bLhCK1Ndi/codUYE
YstLZfv7XzoSa+8HuAzr3fdLxAs6ceVHihtwxs34DHHI2m6Q3eezsipVnygTc4J9VOXc5BXEfGJp
V9m6XzeaTSSrxJ0rnKUJxwGr0WcmzFEsuGJirjaHV9zVbtv2KUluITYkV3RxbYTChQR4XdWeAb6k
6ytKUfLEcn176S2Bh51fU7iXQ6ZlyxhkR0cr9zEzyMd2wcU8DZ22syqe1pg3Df/lFhTigaYLJbOg
LG1Q/P96GkRR2LP02i3tgxkquDyt3T92s0enls6pYMtXAWiP55dh6R1fJgYa5Z17rOpYGRLmef81
okHzAxVAXCEzHBO0JZ2HutAGL2uBPbPjJFZD64cTG1P6zD7gJ1lTb/jfg1ulj936aoluEHy66aJi
uCucgrqZyo74RTwyCjApabhIKNeoksXOcqXSFIfgpsR6P6/6YJuSTeJTOnscckJ1KtC6i+ZQT49G
oCnbPu2qTr1m/XfHkTY9dyZSu1VyOQsai+Inv8THXk/DJWk4bkGaVq6Ws08ojy3wK/ZTmhpXCgLe
jjZlDrWOvu0A3N6460V2So5t1qASlY5A5RkRIdus/KU8s2CijRiESYxFF3ZTDSK3T5MCM/eRUoDI
OfrTmF8M/DFFllKDJnG7YphMH8XN1RfVXYS4XJkIPsbck4hl7Mzcc9mPa5NOUnx9k2zNTcuneQNF
Q0x1VFco2Ma+m176YP/KRvbONrVCOCIqIZI6GJMSW681z1ckoG1wBESnCBfcwucdUYHoZ0s06dT+
cCgADZojBitnlK3tJY9HC/siR8l+jEr0dRC4wgY+lYFCvU3zlG6wdmF31FbusJeQ04RExDGCabui
lcHtOUECP8O8jFt+58uMSrIngps1mqvhBz+rt+U7uQQh5HJwEHNiUorCWTO+9KHBEs1UzbeACERK
YObegw6Q3x2fa7NglscULxxoefbgTOhWBv+A1UsqWgH/3VmxgVRO7jIVbR1E45H/csjEvafTELeF
clXQHhq5uiTYZA6OVbNmT5vU3wzm6KXHyifKY0k84FyoZNvdo6KiEdedTF0qeKPQs+8wkKud/mL/
m45/Fm4CGHMYKaNp6YhDZU/aOAWoyrvg10MS2cQlRJZ3FjjguWspZQGI/tDfLNml1PV8VcNpIYz9
KrCGZdyUOcME3uEoPKlp/5xlQFMajFm/WFj6jj00EkINIUN9sdpVd7zcXIFRJt6M53gQTf/TWQik
Z7DSV7gFixrwhKBzFfc0HrAEkp50MLvsjO2y5dBsHWwfwEFvVQY82enhb9BcQf7GdWuKf3Mx5MXC
OBbZKPMqczz+X+yz3PmcTsMIUDsFlgSzwq1Upy4UYtK9YAgdlsL6hcUdjfuvYybCQ5aRappO9+m7
wynhmY8eJR9UMTsM7iTjrthjTKHEwPD8bDvSgcjhKlFyj+EnamMxKAq8tz4a3/DAcwgphZn2z0Ye
OndqKvIO63e9QKri3cOouOHs6uy3zamB0LOGw8k7ampKzTfsG52Pw8YsoeaeLxDJb7mib2YLhtxI
HG83aLSf4iy1g4/5TyCiafn8E8cuz7NRu6HXyWSpm6ir1MUthNb8wS3/NzQoNctKf0XfyG8jcoMh
XDkRuggipmMcOTOCFUBuFnx097tSbPXAxtQ2oMDaa9yLhQt5+TwQxIYhuRsC/jQ+UBVBg2oVVhTq
2b+5A8A4W5fBOnLpRaiWjc3pD+a/e7bEZMwySkfgwhbT6RBVeerqcJdGov1sIHORT0Kveg8dFYm1
MRusvQJR6J5+N//qplhPD4DzsTbdwEsnmtFjz/AwM+GP87Od8gBbtvdxjbOnzZTgSORksmYoTFXf
DRCDgdmdxyNiwG+GfFI/OqE04vA4SkOkidRr6h0l1RyCsDvHxgbUy59/Exc3XyDImdVGcYXvjkif
DLcSyIbVYteZlt6Ihv0Qukazz6QRukTR5VkFIajV5CYvsSQeAo3GLPe7+1eU2rgp3h1qDM7XNpzP
BaYiYXICqMurGm4m2I561qeeXivHnpQO78W0gIbMnpzDgF/BSm7XbVcHA9TcdCDjFu3mmJ1AwuKq
Ip11VRjDMM2fSxrd9vSPICI2IYDwnyxYMgBkXzD/tcyRzk61fI+N2MLUlvyKOrXs0M9HWRECwMcJ
oq/R7PNN1sXB/ozUQw8IgEiHCUs2pn0v1WNgTI9jeRf2nVJmaZIaCTP3GXEM5mQb31kxH37GkG/J
4CvP5mP65Rv7y9+3moXbVwPqHcYxhUtBE6gD5h0pyh6Hw+B2o8hLfun99XNjjleOpz2AbEJ4zXOE
KyIkICx4AvbJep/XTItAPV3lFygdH+siWyKEygKfoxxyBTgznmAsTSP6QuCRQcDeJrPehZfnb4Nk
sbf9kXFTcImeTBd/+wPpAh2YOEMbCni3uxButlFZ2VOUrPzjipBTHT2iQC/eQj2j4WsBzsWEUbXf
5r+ZroKzOypZhpbvf+2JeGQofhXxQ19MwWNBDA9jwv5fU2JPvNjfRioCOyaXgn+wEJokem1eE18v
r9lEBLRwMwIYa8RXsDJDfMzxa3sSFc9GGb/eojrv4SP4+BauAuf7QqXab0OR18EaCMvvCRRHZcvW
rsacgGBf6nxrGHCFFEvP44sFJY/JyftxjfKuXlD3sjENNKdv5iO/WZsmv3+uy1kRJBR8qZ1mlGI2
QKuz8Z3+/w1mbQK+2HxJXmgBozz1GbiNguto843QtwiQwiomU/NQ6tjfz+lzNDq24sTPUpX76WEs
hnfVNTB1F+2tibg3P29MrvRCiVgd6CjLRdUA+/8Pg+Lx1j9Zt1nS0lmXRjBXOeSJZ86d3rNxy6af
9vaGSThPBSIkVV6SyPCa6WBkhOxE8fxGyvIE2kuBURNaL4PDeVH0AqMZZtwIg1vxEgMgwdJK+svs
eRer2+fnG3+VQvo6B3uE0HhwHhpvoH0OqX0odcJIGFn/Y5yi6Dq9Ajqh0BnlAkPetlM954SYG5uK
oVQM9z7+LZZQpRARawQLtNimHPLVN1FM6PRQG07eCKK/9U6jw/tHusyyo1I1qywsEzCz3vFAnxPh
33TH7CXtkQfj2Vd72hLsUV2TuELrXvIPXpkZZUjQoPVl8L2MN8tnQc2GOUO4HjY6TkgecwhJ3IsB
TY6eWaFMlMB3980jRsJzBXYr6Af/ART4B/6k9Hc+sGTLr+tBJ/URuR3+mO191ETNoa6ye7wwkLQy
mb0U9qHXdbsUwmBT+QEj8Bw2PfxwjCqmEoEvZWbsIX3MLkeiSNCZJpL8cw9gDFLY4d83rpUQ15cl
SzqXrnxkRb6Gy/nV65/5jPLJYX25ZgCv0DKzs4V/cfUeqiNRD6H0O9Qsun/5/Zy6E3/AYHGB9niw
A2pmkTsfnneRlQiRocPEwQgGZb6yXYHnnR7BkQmklUo7DVl5Ih8uIoCf1UnEZHS5THplKgjSRXjV
nDuy1GKGIg3SeQTUxIM1DXKqZcXiDqKaiSbbBFD0Ukiyd/OSxpsazCT4ym9/UwA6W2dhY1SJZns3
vFy/dleAaIZWWKgLlBIqnm/2vS4LSPQYzhPi/vLNjYFgs+fNLW4UVipVn9+cDMfUL0vvAVK9dLbS
eK8WjWM+OiKdQHyaKq7x2RMiwXZFKEp47LMjEdQStigiD8Zps1DimGb4Kqa+vTqJhBbrjQwlH7RO
54/7A8i5OWa0H2c5N+LDG5qNGYufWvktUxxhAThcXPHVeWHbMbEw2dgLjVl3uDBWmYiJ513IoS7m
IacRtoq5+HDQ8JblDAqvYsRh9JktP2Cg1r5iuVS0EGD4EomDmctKtqOxnhDN6K8NAp8Pn6pXnzB+
kefSjvCo7Y/kmEfEXJ3TS3Pee7TM4WDEM+28fJ7mTb8TxzFawWtwK+WH4qM+XTk9cIZCXYdxY4dN
DvHXl70OC3lHjEGlHCLoJyQRMoYz2uJiftVUvcajT/9dvuMB2Lwj7p8n6+9N8AJbr+Mr6HoLKAdw
DDgefXMu6huiZyd/N3Ck12xCgHFdUDxicQwANE6ParPcHcz3RKHhbPNJuUAZuP+hGKvluWZYBfkd
pR1yP+dGMu+2JQlKSTaA6SwIgKf9sMlYrG0lQdH5f4PSJ8FUz38syZhBVIV0IckwYEyLL3byrAXI
jZQmULkNcFVSWdq41Qup8MT9z+yz5HXmppkoTAu/KNDX7AfOGu0N2BqliMSABga9jSOdDED0HmUH
bKx/wbKPbwmQWJ0pZinVxYOhSwlsrj/2OacWmpFZhSa+d8Y0P1MtgCrcKvRXwAodZdR119zJycG2
DorGJS3HJw0cZgJi4DiqAiMLrLUkOVonBWh0o8i48pK5T5bgD4dy5ETPMRmD238v++dFy0uFnK+2
`protect end_protected
