`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nwI9apodsxWnt8/qZ84l2L5r2ru1rYRvzH+cIiU2LZ7ZFrYGVhrKUku8GacxvPmk04mNLHGAUf3D
0KN1yrZ0UA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Sm1hR/bXnEX5hSLJC+m0q+qTo+GE1jW/bGh9GYODVR1B61WO0x3DI91rmMkLB3jXabqZYmZaVRnk
N8AiDf+w3tD5cTm9k3UfnHfkmqEgj8LBJAWCYHciLWzjmW7DKTQG5Copg5YaoAmLrkH/R11p2QBq
US3uTE+2f5z8QlQwimE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
y/EngzI5VWuiEHV+TKhmZG2qH1QkzhsLqS3InhpMlNY6l/FsFenjJYgIcwfRB5cHNIe7FLSQt6Ne
y3HMmpsqF6xetN1AMKtt7yIa7k99d/5TC5vyU4dMYs9g27cqHYJzk93esgZCvjIZLHpcXw/tu9/b
4U5FbTjst4GUWQQ7e+FOVWa1BC4H7jo6ZOE8mZ1oMeTUDMRBFFBQWv4xUZFg+dKul2euXKFScShR
h6tknaycBcdNbA+6dQJo+VgrTTewvfrkpNyifPBwk9vIitRhFkJJJVGsR6T+AF/UJfY5dEYYFuu5
J288ggKjbjEUNQnIyNWOpZiuhpClTTay3laNkw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
htKUMvAlzdN4BbAAeNmEM6Yr1UUCORwvd6+1cV737AnX/e5QyMGFY1ZuaVzrrzfIKK+VWd/bFDYR
WeL3jKvGUsyl0cMQ9jcxLrsCI3RnUD8yDbbqyDu9KMj34D7UA/k879CbEg7mJQsE/OUuwmk5Rusa
S2E+UVp+HrYNnNymuLmmn6wOTCKRZjZEMW81xyRvJrDTTqf12SjMprM/ubdETBwwiEzoIwLeibWv
EE77NEiYVwYpzXElBkB+JN+riXCrervjpMbAzHbeomW24pwXmffMMvkj1nRzaEI2QRT19Hpc4iqq
tT7PSLFxC6iyyFn2bd5a57kSCEK5ZaaxszxEVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ST+OORnrF+3QguD7AuqTgC907V9FPxT3xpP2TfPbwAQB2+m85/czQ7xrlMYLNRNl2qldRPC2JAtf
yRLJmvKEgyRtR6tv/9gg66CdnvMVGbBmprZnmsgKpHGXcIGIVm6FR+ifL/5pZcFZyTQCKYlbE6bz
YNrIQ8EskAk5YXNHRZU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Zz8HkbKk2BMn9pYqHdEWEMFHnKjJed8tZnBzajqsks1G6q0CzbV0FSYoWS1nKj84tIU1JkBaGDIt
9sdF4TFidxOJyhtrmpNfTChKxpMr41K8vo0yCOwdi29v/VShuI/rkIBCSgrdlmTBWBEgiBS9aabp
Jqqjo1ol263k6jlcp9rOjaoU+lcQMEXCkHoZu/V2+VWtTqhoSiWKgDQ0jJptGQig3wemEM16ctGQ
xX4urrzlEYCVTlr9g3mn6x8NgAjEFjJqmg1uE21AWGXfsNowkj2dYZLCXuVTF108ULXlOgx8TBHk
tPYc56T7eylPXV3Y05Z7agtvOLTYldGNSnm7qQ==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VHzNHo3jyVixjpbjlcbNuO7IrIjCuYoXTAjRb06/SIYnbUS1pXATLQwryf5S2ETq0CYvThlIAGS0
xbNOLpEIhHMaY4VNrUdhUPBHXcXHWUCHudYKaUCB/Pk28QZKLuHYt3FqZh6wdzI6AFJdP/pykVJb
M/Pyyc+uLtqsAqyWqtJ0puNrBSpFPSM5259v7Gum4dwYGluRNUyJPq0CnQOQDcjaKw42cmf2DAtX
CSJb79mvoLdsFiW5ePQbcfrrcT/FhIkNj4/DqMVl2EB85zQgcPJw5Up3lLGw0Qd2Cd1jeq3A4qcf
LraHhfdfhy6tS33yDqFUeXlzvLfkicvxivScIw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2020_08", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ir7vg+6icGbLB3CLLO2WEVH7p5OyaYzRs27g9ktjlLGEA8UZWJVD/LEebYJEdrotzhB8SWmHZMDV
/tU66bmEBeBvDhzPDFffP8JEne90WI2d4WsOz8gc/qUmQrWkWWpKaGeRzRKobk6HEaC+nXg3PqfM
0b03fbE0S205+4xE/rEnuHBIRBfZd3xmeVaB0HKBt0SGPD5SSQQZpPD38QOtCELjuuuA4RtmpS90
kaKEHc7Je6wpd85YQOJtbSfSfwms8QmBrV2vuYX5vgvFoWdrKhFu6ei5xOtYRK3gX3JKdEXLebbV
49uISo0iQ96Wfdc+51UDQD4Z2sSmPF/BKuQ5nQ==

`protect key_keyowner = "Metrics Technologies Inc.", key_keyname = "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
LpdRmMYH4gdKs52wqPlK6TsP8t36Rz9etYG+uFXIxoYPOw77GvCpHTnPEq4wgKvtHfjSBYM58T8o
VFR+rx+dgG80Vv61h2/ALXu7WMVNRnj432YN7jUfiNGlmdGjYf7j5bb6jDSZd9SGg9hOG322ua8w
FL0iNhZ1+8bqOC5DHZhVoYhtH7wentMTqEBB4I+Xy3zK2H07hbY20A+hZ5iviyCzHMtmQ5LCJzAb
8LeBnGRdOv8ntIJz3n1voQKFpamiYGRWqDwIHC+A3vf0VlEiw8M53hPC9SjoIQqQxSnkzTditbkH
fDStRcfPfMIOJ9yoREe7QoWlh0XCwpflnMvnNg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
lG1UHUIfxtobOdZD+rmMiYrCMNEN9o07Ksv5hjN/5LnCctJu6Yg4/dYybj0CFSQCoECYoy87WhRs
uXCay/u+i1BHK8AihSkKDcYPpvAFzBShXjpu9bdiHWOXHkXvP1ZrDhyEcgNPZje+p9xXJ7cmVg1M
C5QP2t5GBMjnyXTlOh0LgX93Q+b9hpJtbUoGV/g1kAG0OIvmAAJKzhne0VvZuhG7fw/l7dUCl9ZA
/deMMhPLmPmq+yuwMKuDimVOhzjLuJxAvXBfJRFLmC6RoSBfYW8eQTbdt/5sG8uvJqpJ2EjfbCWT
o6/cjy5CQwLZjs8FjXXkQ2u8OVWQ099JFl9QupmdRiYcmeG2V2qHEB4jN2A65IiePfMnrEFtH9HI
ocgkbs+2w67+SYKlKwwlvxtGyX/NMjSXPG3layaRewX98LrQ4cysJ35KFoVlWxNpf6EiTCJjOECU
NprIpu162EL1aZvxHFGVJR5U0wfVF6gdlQ37379QCOkdf928d0vK/KsywC/anK3zdcBIVBg6N2hf
9FwY/BErTrcojqFmEHFQWV4jXHljPv35ox98FptqJqHQT7NRnzvwq1LP85jRCRApfYjU2wtDlOzq
/jAS2H5Eri/UJFkyrjjd4qFyaphyZ/dXSsb3+KXgGsoQYcr8irKhbJk62G0SLAP3sFTgXIyKVmhN
asQDeCpclK/VMkFVwoWoMg/bZmVv0CXkCrRY1UCoO00wm8qd29oeSP6TMByMEJhRJHiEaTVKCfTl
wtQ8YekHQC5OVFrViEzM299Agqx3Dov98Fvw9QYUOEjn+swcmkpd1SYw9xFHjZl4cYfuAFMe7nuv
VNYyH9br4T3t8KSLRr6bHtIvVB7hmKoSJQhdiVEOo7jTxAM9q+upbjPdO//8RC62do6idv4YybcS
nMTaO/I1pKECs1CBJynhIVWUpZNvGy2z7OIbJd6tK2XgKSXIlGmXaEf6JXnDGaZ4DUx/0o/CMuG8
3EgoDks86RkGcs2BN0Dmfe5yXAlV+Qes1e1GPZjnTTpBpRhW3z0BI6hQFBg+ofyw76mA8n/MAye0
KnXp0VMQYr1wQEU1fO6sIgCeIdpId4dTVNocNf7XTEQBZJKpGpegyV7wCBWC8SiS/O23nZpJKVg5
jnqtPJL0x33n14OUQnZcuIIYNq2jUZ1OxXmD/7cVClq9Y5nq005vLz6KbBYi66C7SJK1P6qPqVAQ
K6hSIs+Q2Ms3axeK3XP5Cjd4dQboyehAA8NmA5paO0HH21HU//SqL2Y1aDTktyc15cFLn0dAOa/F
MpOmVWn7s0hCyRLof23DwxWNQkqXN6HoIZOERU1H3kc32sRnuRG/ICUyiI4dk0aR+Hno6K26xYGU
jve5ynlofslY3iE1mMrnvjZ9idnj5A1vu+eJHWA7yZhfhtXapfAN8UaohNwswiU4wy3AjO1P+Ir/
zh5oEPUGeIbJBdX8PQep2XPNO4KdxCBWwOb2nndphRdhE/0bmrAGRujCYfaE/PcpgyJ9evNJTLdQ
paba2v5ukh2nl3NJVr3xIe0/wVVXircwF5fcfwE3uCc3qNnY8RLRev4b+GoLYF64ZM8oUcDddopL
BpT7njdub1DvRZJfnh5bkNoiq5A56hv8lRhzjIS49xGAtEXRMCYOuEqHyqwrtIX0amUf1xNSzSrW
qoneO+dyGiIXSycoxEdp64SRoGL5F6V93Jkg3ZrzerkQQtpLos8/WWTxdus9b9pe1beVJzyXyrjq
oFMZgQ8zBrtqxMqjWy/eWkBRP4wPMLPemr+HGapiIzOoTvfgXMfue+t6DoG9hW87fDdI0KqP9v4c
Q1PINtwx3YtENMfOON3m3XvbD2Kxvir4bfgkLgZQBJKgWCivYMXKzIa0dZS43pzwnpww1vBRddAj
gvDq3MCHOh9c3gtuvgc7gxxjqUmmCQZfCxxxtudwB9TzFL2fN8hyKiOmLSPMuCaSbMKSkrJ1VnBK
zMwbyWpZ3bFHPCg+mOa3ccFopO3B3Rb+8FgqZ5Tm7pqJsnG9+ttPneOnqkQGldqhwDMYonRi4fFW
q6XG2sgTAP7iTENvVc+b6mtLwb2H55omaU13czseSdBUG9LuuKRpT7GZwJhkgqf1nzYe6OlH5g3d
Rhe3rz0raAlry3wDyb7vTbhYc6kGz4YUy4toGV5F7Zi455mPHffGPx4OUdsUVPpW9pAACg4NhcA9
S9Z97ZJAXi3EthuGj/3zevCwtyAxNrG6l7GRbY3LFCTppN3B7LmjpuYTdar1aIr9iaeonpqtUMnr
9rcU/s3HeFgCal6v9fq5/HAmMQ7D8eFwHPGjO6o3v5iB9ah33W5lqS6WE0CLOGtWG5D2q/qYoC5c
z3dgo84069uktzn/H8C/zBr/a0Euy/rNy6BEmfF4YMpKUXTd6alietCcXyG3rikyra2FZapv+E/6
Kp5URXhfV+ZcXgBiQc99AGKz52cwGHt5MNgecd4bMZb8Noq5GMKMLnAyZQZKQ8ztDhjqkNHRl/N4
DFpFetxPARvNb7N1YJGinzV2pXgRDLJYoA9QLmOeUg7fjwY0UcKbbbi3aF20K2eMtlRPw3YojVPK
Qhf/iYj78KMnRhP6awecYFL3xJmm13zt4Ip9yeh+ViIRhqrSai5Zna+JF6UbE/fRC7xhXmtcl2Xk
2V7GLjs6eupTCCiOPNjGF6LyZq8A/wgalV++q3QJTFJqg5ta7pYB9agHOJ0+AiPWOxtiwrYfTUNg
QYwPxaOScsJzlnZ9gQwyRuq7Owpckb37aLApWVe13gGK6DHK3pjwHiQw5b1bjGetGV0jjsRus0YX
NPJF+VR449jn5hbWgLlYjnoidCk5TjaQz0b9xA36lDRIa1DId2Xd6TLsITlpkdtO6IZUMwkM0fUQ
q+DZvDKlz+lmnbzRpdXVHtsDYcLvrEp9idKh7QiVurRfPI+u9ALTcRnHkW4q+svIP0PO99AKWJqZ
nIRghA/mc8PHdU8CHygwM3Fa2t/7Y3alrYc95vuEAYXwWt9F3vSGmkm0E3D4N2YEEU1dMWVIdCOR
yuIYA8Au4Vf4gsLrTygn2/CIe9S4XUopvTCjR5cJqHGK4dtQTBili5kLTnFZ61b9Lv95c+JmjbJq
Y0iy1S/ZQfDeP1VzipO0UEQAnWYDclh1lcM4xc4fUCdF1gOeKtQK4GzG68hAILj3TEOcRoibACnK
oEzim5GZjbJCsRF92g7zDrZiZv2mr1PHmZg/OVriRsCcM1XdpjMcJsuuSsHRrlNm6KilYQigvwtJ
6SB8CyzEHe5Hv9AINB+Sks+ALQIOXWM4OQ5RCAUrs2atnTv4aFN0el9s54J3gx/UrkOCs3elWGep
0CFy7RuBOd5fAzMjCno0pWQO9RrhCPQwankve/pj0Q7LauimPMGt3dkFuY/GTsi5pzu7T/Ej+SRR
D7pBWfxPAKrIrbK2z62mTin0XZPqBwPzNXflNtgrHx96TMp3YEnIfbN3IKhSHly2yANt8MJqDDFw
u65jQwP27jZOQVoZkVVZxW7unMnTvJFRPhjsy2itzPYr92kCXC9zeLGFp4y/o5PrwjAAz3gf5nQh
cmt8gwQutoFsBW3wYUUrZwpQVxtLxD3A0jB2S5YOxL1l/TJXNhErsQ46M3s2P9Cw2O01jH1IEIIK
gJRd7QMrU//U7YOGOEGiDT25Vl/TnpO09DEqjrGtwA7WzH+31Tz1DW3gaU08Bjta/GOQYPT6Ug07
4Xp42Mpw+ItVYhRfAu2KBmy4n9mocvv3cvX5zIHy2oydyf1UCKsirsyzI8IuridKioSBNqVgsLys
+T87GezHl3k2Ab76h+JQ/ALRkpgEWii+GZUIUB/JIOd9ZB3Gz0bVSnEsekXx5A/LBUSFy80Z+MTa
FMyGslP0tPEQMXwZecA7pOSO3HjTh3F4vKlqUIp/yovOXSEqZXgedXq157E5QN0hWy+UuHeuGjBC
zMOejdP5sqEZfRtoh4n82Zqz8t9ZZ4OR3VWSApsMc+JkHfZQ7wK97/pcvpS7C7+cSpB/Y1OTr5HR
qyJjUQiMFffRcf8LnFDrf9UazNMHRc8XKxu/1rGf3Bhy5X0tleFYhv5ZUo6X/67iKXuvHgUoqqdD
nydiZXydPOZ4SvMl0y8WZN+0vgmnBljYJp4Bh2Xd8xezdoE+bEDuVKOUE60RXshfJik+C0I+lHp/
B6sT73+ZXYWFDD4orTBwUXGbm13DTM7hVGlsBnBYla2ulKo0UNntAzqW/W/sJ29+yR210W9K/y/K
XlDdClMXQEUP1Wmu7Kq+JeU3icjuJQJ954HmU+n6kgnuf0HRcLitXePNdEFcNDkayflKY4T6l4Za
tCPZM8tYNtdPsnYd4c948u2tXY7chmBk5R76FQ0Wjo05VFjGvp8Dbzx9QLq0KzUN6kAwI9ReD4TK
nrij0AeDD9SabWC+o3e7QlpCuMOcRzwbfhSLkcYYXgBL1+VKk9R3Mk2tT98wVw5X3k6wEhK2Lfxz
cM0RmlcVSNmg5omfE/2UIk+aOxah/rdGKCL2p1mdaqWp6b0sZHx09qc9Qri4ufQdM2qHitByFXwj
vbhvUoCvaBmFyBWXdynDgyCkK6ZmZxxbORiSeVCIRIC1apv4ECsHsTdQyqYQHcaSdc5xXkGBa3Bh
t/4iHTs0L2JQnfXhcbN29WtZsj/JCUIf9mLoCeRzXG06m4/2YpjiS0B4KlCuWC1++bUDZOY5TrGQ
iMT6bfFuJVzw8D58MY3Y3pimYjb6YJlAvnd93WQZIIcy516YYf9kR0sXr1e/PRPAlWQHcwJLyPGN
qR2MFwUbUuVHXQ1aPhHFRlyq29UtXEXxLsuM4yzlxF5vWhisaBx8FKZVGvxgTFYhu2gGVYMQliGa
fvd3BccjT0ePnRs3nj3yJwwS5HVC2lvi26OqRGEd0hlBYXwA+bhaSt4hNitOJlZajVaZPyuY8DP1
twqswtqcQYYXX0nSfVScR7bROKzPoXheLYuZk0GyWwXRIqsfhdiRZOq0OiPkjt+AE2vvQ1xxQ+2u
E/4jxfJ58CFqD271UbwC+6QtOAfAXBB+otuZSdXBPFZh7A3Fxjbl4gWRVwW8xabuqv3dE5cB4z/D
+x+NKs4q4tB/SIocVluyVYg+uU28E7KOhIk007JJNVdty+RqWRdNS4eS0VdscUq8XJLUSbw5YeGL
s3Dhh7qdiBq3BVHrrnqjcZFOclfSC/4hiiYgkMdrOKrg91Av+h5TNMSEVt5kdqwMvcIHP8LRgLAU
otgqVo3LpeLW7CGvHnFEF+tetLKbxcmDQap0LQCvm9/bNY2clhkU4JoQXqJ7jaYGapbA1GnGOwN9
HCEfIVgxKLEO+R9La2r1LfDm+guO9WvJr+lbXHxxV+W2RGysuhIqdHVAB6q+5iP0DHSgUSwpgB98
9iAp/lfg4YGJpFbeBjiGAgT6CShVTfxJ9GZeUl25437Kc3AXRsJReMYRSBUZqlV6jZNK9zgAbTN7
7ikOGI/LYbzCtufsDHWm40vYUtJN67Qvkb/LPlEXLaC8sAtmhAeB/gsdyxPW3aropM/cVTA9yGxP
7ek9LDAXzjbb5MPVf7iAQa2Px2B6eFNwtdmxg6v51iDMccn5lNnhavQhSPlYA2fJTMzQ7IwXpJfv
/eLb3okyjq43IU/0vL9NfjNeEvyrx/tGXDacu2LYOhR+gfth2gUy/gWvk76TZqAco/JNqY3dYUez
xp82VQm3mrKXi1xuuuUWysNkzsq5Ud9dQyYjrc8ks97u7NYmmyWGOuENuKKn0a4jLz42D2HqsLwa
kh7YfT7biM1IVo+gO4Fbu8U+B4S42/QyCR57jc7sjPyRvCX1ubyiDZyk99DDrG5oo/bt6D42tOMs
ycA5RfszeLb31ab+R00iIVLe35OouW+QFuiI4fbnTbZMovMmwUPisR9bNh/ELWCmAPfPBcitlk9c
zIMmSBrDW3tQjm0O/EJtaWMEDpkP768Nm/C/s9cTEom7JTa7l156a1s7b8Cxlm6OOJsgazqdOsWj
u+XN2wuHfqrzx3pybaUtlL5Ie90YN2jfaPx9F60HAJ/gKAG1BOzU9HVBe8zAYdIptuh0BhfvFKMc
uvp3LhPcTtkDPFxjYZkYCgSEjnY+QF44Qg0WgkVNags0+QPoUgjpY4UVx0+CCDx/A4CKMqQ1gkgX
Q/1//DXjATy8zlkXUw7jsHP8kxqHEtCSYoOfTgK1nsoaeoWnMmTyebgq/XiHIRxmZPW8eeODi5jB
eu7euDYc/AIaDaVMkze2a5YQhyCEX6KujW0Mxh9WccvMAimqphfJTX0tyFWmS3ftsJDzjXskeXud
DzguOj/bedFumFFnxRzrffi64XZ/nIyeDtxQX1zm85IZC2Nomio1zaGq0aKQpnGHTmSdxapR+fei
IfshNVu+B2v1gbiicK0lFY1yI3GzWTwDZilQc3TU/6z43gN/xQK7TGw3ZQ1brkTJbwb7zGGGXSWd
jZXywn3SFuuhtjE0opjrSyaehfeUPt/Muq6/eKddKiWBWPpfbJEGGPcLlGdJle634fq897M9L0Yx
zYfE2cAUBgOe47LD7ul2y+1FXY2+Z+QSBT/GPXOHdxhpVwJfshQbqwQXqqsL/ODPXF9jbmu3Oh9i
8SU65Tp3WYaiaMSOw6xLtFdrDWHjTnI3+5JT+i0BpqOu2ubGGe1pOCsLWVbrQa0OaLkk7cBF++nu
Kfn9s0/tUItAbwFP4kZe/oWLBYuAGiF8NVUxVFlJDh9MazwzJRPr5m+frAZG93pAwk2ne+olSRcc
xkROb1sx57LmqNa79XKSai970mDCbHgNuVBDAfbQJNlSrUKBtSg4K/zlDxDVrFwt3rNqZZKctuwe
Oi2jkPuk0zQbV6dNtoH8pos2jTIqZB9w2KoymgMoNvomRCAiNkwT9rgraWD1bpDPOZIjZmI7rleu
H2CsZ4sROkcgnPUX1f3x6CunJhBRi5iHMl52E+Yr+NlcsB8Tti/XjI9td1kJQSZVCSmbeKp4ca1T
JNDjuhXsrUI+3kr7OJK4nXFmijaeEOqSPYUj06bNbIH5t8oRDP4zX2+y1FEqQl9DRt428shgxmpo
ywABYTjM6Ez9GZuQS6+F0E/5ACfHZwT8cG9yEyEIlehr1IUXGi13KnbUr1vbn6HksAOdVerwX6Cv
Pvb28DlBbILhz1Ba/2tcjM5eRosYGyZRifV6UgpFaE39irx36ltZaHPU7Jq1TwQ/yx0CKJfhfSSu
tTIX+Si5UlYujmU1kWXuGufPdimf0KNJDpNGR9IpkqP0arvW2e4rqbyHZsMtTrew8yULFaQ6fRB+
5kf0fMEx3fWxyPSztl6VPW6ItFrlHS2JIjAYQ5KOg9FWSCwQ3q6J93zKU9xV6rY4u0o4gEraGa8V
M2GiUrkjU9Muk6T9TzEHmINwf7BPdgV4dVxf+SiIpuw410Bdbi6DaKNOZbzU8L0PKvGuhCd+IqH9
T4p1ICsks7sqTpUP4/UUNj83igqYdhMVrIMz7PfsBHs/G5q0w6jXct94h9lB/Wyhqb9QAjN5Y7Jv
gmCxVCBwN0HxV16rGc1Hs0lXg8A9BOzw4Tt+jPraQka7c2QoxHGAZtkAU0aqzDUwgximF2BnhPrl
fHoY9IgufJjrGnoJTRM8MOAB9PkRKHnRV923BXx585e8BnN/RA0miP8qpmMKg5guywM0HYXFwbtz
GjU1s0Cek7ti8h3mEUTEo2WIgWlTlCjz+Lfe6mCxtRq+4di1IORRVlCnYP3At5Ty/3OhQE1Jz19T
/gSJQcRCZGjMTSQU//5zZN+w303bEQxfR3aYfQWDRh6liFp5ChNyiLTLRScXt+ruC1GwHe/fVNJ8
0E4qKJuqXBZKqeG/peVMRw7hg/UGA2uP5hDDYDU/b+r+lSpPw51PLz+8srR4ZDehDDaOTNUJG1L1
l2eJDuozD9lW3n2DfvmqZfxRnBmv+qtAZrLTGwWk6nyb0iCHW2hPmXm0ivxWY+fZ73dHHHL+YbE+
Yd3yQ4PjHu2IHRCnH6ief3SPXLCsfePRAUuMADJiPo6FO6zm3rhSaZCja2NqzwqUZimzg14AhY03
UdtdaAJaIdZPzJDUhamL26DM2omTSGAh6mz6KRuPc+e4FHLbOY5mtESGONoPHoe/58TkoVOdw1Ye
zYnJswFd1GBz8r5K/30EJLuiGjXmBC3tqBGi6kZQuIZACHFLCzFYibqtcT1h7AFhmsQ4aW7R9jiU
OIKbQGSR2rBWl93DxHywfTN1M3okL4V7tggKboZ/CmDngbvLJUtX4Jsgrt/ZRWxvGAKwKUf3N8Q7
k5yMdr1SMVRxNxFp+lpXYXvSX8BlPltE5Jso97Dz1AkeLNb2Q2zVijH5+rnv2fxtgtip2xB2GwH3
uTtdqntPKmdYBsmMI+6lLx2NT5IgDYsQm5c4LWzX9K3EBWM+CJZBDm8/gkY0CwCk2qeIB2mLZQ4H
gQZuYmvZmZWSnC8SGKQd+1EhG97MK8y9rBbcQTU37soGfEKsTf8dTRRSLK9enLth1djDHbkttLWq
2DupDLLtJdbyXYeVVQQxlqzxknxeupEcB0+wYIKPQ2OVjMgvM/gnPDRW0iFNnI4ISFdDV1cPuo6x
G0gC003pYjrjQiZb6t7MS/60t1qcDsP85C5syk9RpsOufNWoKr1noauw56giMCu6rCHKxbQWyxpe
JtOBsTQO2aW1fjKAl5J78Nc1jOZpE0ir6niTApn1Mzbv7Y9IXZr/CAJEtIkafOye9l/GEg2fSxAG
ozTP50K4u9VmjuMkuxLYAmYysW8fjHE5Ms2fEIfnIlqLnZM/eHEhBvuvujQBeI+g2xwL4VmvKMMf
UowywzV0LlWet2x4hn7XIx/KViZOk6gini7EfGKwpIqJWl4Yk6ePD7RqHcMuNkJqadvPDk8w8ZKL
BI9EY4dS9AWY6tQ9rbIlvYbXlA3y3SZz9ttilEGvCb/aY/aOC6JkbtmN1UAjhTIL7N0cKkwyhWpS
6HRWbZYmYZwP/aItpye8w37YGwhkyZWZJ6JKipycP9p0u+ApDUs0xmcPi4cNi4aEe9/1n2cdMEnw
jJ1DhB1oLSzxbzmGqz8EbwCG/CbNjjkkldEJUaOTvHds/21s34H09Yyp8hO5pMEap+cl+CHPkMmQ
insMyYIwdzhGxOo2XcbIkFSs3XVytiOmRWKp3FxoXaus50tslJBa9x2FfZKlyWTPHqyCwoI/wMFr
H4QDxa9o9VjCeOLIn+4JF8lrhKoQ/X42KmSP2G0uDZIKx3gATLLXg7CwTs7h46kFGwqdZqlB3Om+
DB3XxlWFC1G1WocyE/nZYpUVC0YRkwJC0yP/AY8e7drCkd5NP8tuMYIFNTnPQYp6JrVCMb2HxyRl
xT0lvQ3nw1t4yXE3CfhqZCywbWXDws32Be+q9l63+oDTLs8hyYYXkP0txzWBYdldO00y60mSb2AI
4j8MkomHPZ21s+Ff46Wid7vJsWbxwxUxBLKq7Rv0wEz3rzgXE3eh/O3B6IY+rDC8JoF6EbGquqHy
pxtLq3o1rg77Y0RkvrxNdOh6Bep9py7VW8+XzyjrXCOP03zOCcy9etNFU1v02E/rOMOU0WqwhH7v
Myx31Duo8zOzQE8pLskb55YpBMr4WAtZFbXI5ZlrhaSH7jSX/sumEi3EHJkctJlnSK4RxSkmnYjK
gUZ3kGUaR613NDv0/l7tVIw4YAt+k+cg56RfKdUKiU2ru142adUl1xcGl5AAS3ovXUOZAIB3GDyR
hVEEhZere3IU3SeqzpCX1Ob3ZO5xWxkn6xPeU+29NbD2CUzd3nKYSIw5GyebiNgL+9LKND13+2/p
91aQPFGSGfhoEQPS24V0c/SqXY76FjoxkPtzxSZP3yS+E6Cvec3UieqwTPKvemWkdAJtPyyFSeGN
JaBK+dS5hrYB4b30+5XDf7Sl/+e0KVHHEiSbtmIt4Xn8FhlCCt2AnXmE3vhd3gQ2SboEod/I4Ed1
Uji9LIO7iDRUrMW0c6+Vh/gzvRfO7I9LCXtWVWydB+BrqltY+WqC8dluE5yiw/QWVeHdtKXLK1ns
hwSl+vt6JqSydjFb8QW/rNsxP9f0Pn9wPBL5bxnAf9vlxJp4Xc+64ovKrmy3gU9COzEUddFFCCv6
WjFK6GF1vKg5mTyJGV2TtEeEV1ucDzOZi0iupxCijzPm33qg/PJME0D8zcBcuo0zEIdfilAfni12
olvQ0TwfZu2DTzv8HJUBb5hyC1ywyKRvfyvKjMKdGzhY6MP/MaCkENLJ/tKZFT73vD2UXvEqf8qn
NvQA+JB68Z+EMQ54Om+aheU4np8sdW9cN3tIGajQ1yo+7cfJqc8d0ebPOsTUAEfvrXNFuhLWCRBM
RSN2FLFgmFcL6K9Zj87EJsKaawsUAbEuO3SXgnp4UQcKnNgsK9J5Mpve3Hq7wPQvGWinSCbtW2iF
GUL5jjrCDmym0cT1U0n1nsqfl9GEzOjX8zBOmh+/3aBcemYb90ZZL0aToJeVKHoQ/Z4ZbXu0xd31
cK6eK08KKNXeqDr0m1duwFjLQJdsInnQhJuMsp/OOXLhKXsDA6SPFyLarIqqXbIeBHwU9JXgb1V6
i1JWGE3XXoEGObcq+HDOp1KGL/aq4U0l6MXR4Q8h81i6fBqQ3vY1JsFqccPsCkMSNGnpMMotVfHh
BTxhMsgGtphJQLfZk2GgNrhabbfazyn5QOG/0XX8K2IjiGZw516Xwoff38pLqCnCrWeczZH8A489
u9X9quGaj07E59WhoUe3hPcu21AMA2dWWbMBmwy5YPPmNJXlOxG+Hv0PfKQf0/hdOh1wm2s6PEH4
T7eonA7LNHpDc9jp6SrPw1K6KXZUCPt/0Y6D+bL3TB29cTYUtoqsPFXJwQS05Nl4/ISNmlqtKUen
j0Bwt8VEFYGgDxegypHBLqRSqNTdVOMU2IgqhzTn91ym3Kfh7qKR6SdgKvVsb/3IPy8q6awz2Pqz
IP4Ff45QLFka1KN78jzZ1BYzFSyS8FST/Mu2KqBBe0/R9movM/pV2uKHs6YQOLT06VpwINQNlMCe
46x9EsKr4N0O5WUjx5bWgpZ+FGYil/59os9MxW0oxQHhpe/zydFD4W5sxMWAhO9hihoayidqPubV
mvtjp5t76HfbERUAO4fB3ynQxzm7kXxtjvo9aCb3TyL4u1NN3eU1aHfJGFuas/3DRra9zGBL6f1+
EqKItUH7VGfPfM0Lqa4XY3g/BZqAGgoFZPtr4RAibKaMoIJLFJBTI0yVuLOytWIIM3x9wEaG/xfe
ZOvB4edRb/3Sa92HKtRWz0oMbejArNh35oJkC4NZUCjp1YQ10gF+JpWuIy4Gby0kb3uRew36tqL6
c7rVHfiwlpAdCM7dFROysXkASoe5LbDae6FxDS5tqPoVwKwfbtf221RqQx43VCIaMPbgnBPWPMR4
74sgw7W9U1EGMUcI/aeTIJfLR/E2va2NzbfDcAz331pcZ7L06tXeV3sbTy0KeTfZij0qp7oiPlS2
FMoRqGtdv6Z/j34F7yZC4MVepWz59kaydBu28rYe4WbKub6P3tfdJPxIXRjTf4rajzBzRUA4sBeD
htcpi/itYOeCOL1w/lv5ICHGya6CCr4dIxIjOZ03YvbOj4JXM+apLdy9kqCmug//3J0Bqd+YjUto
sAh7EQ65D1BcZA924aDQKz7VVVKHUqtfYp8JNsScQYIqhPJpPS5u5Tbe1Y3WWZpACNVE4Uv4n1Sg
JPYPpkyEJUdMThIgVCiMH+klZb7ua2IUNPLCXYMp3t0+DdWLaaLhO7/AavLwcBPM66cSXPJzXEzA
xtl4KLeZFitya/26dRkNK0KzWErPe+FoCp3I1FdaC4gSciXjYVA9/lQNRzafy9oPlccnbXIoqRl7
KTMb3tRVmTgsrkdj4LaENCgQ0OEbluaKbs1k3LvtUf0EFhDarcVrkA2O2Gub9kJUT7QSpaCdAlmS
u6u0CgsIi6oTfUWqvmm6TjUP4ngkpnQSlwqpAdabLrlD7RiQUX7toSxg1TD9lXd/QpQ2OX3c6NK3
uejL23te2XuuEqqnFOlCkh+VeJdpqfNeJMQhhttSxJy7dAee0895BnJG4XPGuWV1WZDSw5Fuhzdg
AZ83Q0z07CX5+3E4dQE7p/3QTKHuMNF84J1BTfehQAg3qeS0CwMHCg/E/QLLKQBH/PJvpuU0vdr+
advm8OXrxYIFU2zFI6omAWQGmdnbTN4F/w//dAPNtHXBLCjU4xQHLWU7k7MgB7tIGR1ucM+CKB6B
suws8j9uPiXM82HYEerRkuH+3lWqaIgCb+McwrMTH1z8O5Dfzoi2MZxFky0BMEItmZkVr0b2ZtaG
wtGWGUnQjEilMqkwHXkyzXBDr75adPwp2nTLbUobtSCjFH3QGZEpQ8SBHYToKsWNQV1qr4nsnvRm
OgBwAVj6jwQVBcGnNzH2GgVjzNE6j5LvJEW3Y4DPUhCbfvz3eKXELKDs+QMaXSqABQQGhBZoM+6U
keGvYVkk8rgLvqmvqv+HuOD8OxkwaCm5DFgealwp/E7sfVkPYV9ryQpOjKJHyeAPnxevLMmZC3QL
3BGi73mMa4vA2ux5OH1UuZuQEN6rfv5A2xzBC405ufgcE/CZqEnIRukLjelDTwjeXo6vBG27arc4
A+fqK3WTOpRWPJBFVyLO0lsvNLV52imm6BB+WReMpVP425pJNWqm1BpN3DD+ioy3VUzE22IR8Bfn
XUQk4bRnIicHYW2G1GAP/d8V0Q4IdChe7DXAGToRcXHMZmZAZ6XAdGrJYgC5TGh01oEkIWqO+BbA
QG9y8Mc/ijtPOXOaJjPfzmfh74KIQaZIWub1iF5x5uBE+ElTTm/rVBLdbQgd9mZ41LZLLPKj1b/F
QiuwGPpA+XyoACmwHcdglNxstM37Lo2PRm9qq7fssDv9QTfJ9RC2reZd+1m+Z7xgDI7rWMoq9XlA
PQIr/SjKeL7Q1PShzAHf3fHzy1i5rSkRlSVxOfpXsaq7lJ7LKDlLR0KScjdo5IQwMr5vM4HLE/F6
/RU16TpJpJSph2Qm1eeUJIvv9fPUBN+sg54I3lQ3KVmlz0KIllY31C9g4JFHSQ5Y42e9gAMCGUvE
FmG0T7m3KqVoDw4wEfvT47RhHwRbQ82OvQgubGpQyqrBl3UOcG2iRgVfwvhmmEcSzm8x8VlPeSvL
QJf36RnTRk27eSIURBrTmWk3y8jkrloQSpNCSPmtpjZYdt6fcpA6N4V8youd4qNOOp80kcQ1svwP
Mg/QF0w9s9+wpavtYlYJ+9ARJhjYqN42pAX+WuTglROGaJU1F2fdVJ59LdVgPMdEk3rrvlSJvo7i
ddSv8W04KtiYV4c0dlKyo3t2ZCMWshidtkIBJaVreJPVP3POsJTa/gZV734HtfHjmDihsYnL2Aq7
1b/WaBzvnQz+SYkS+IpblwZ9v2Z/myLnrZ75I37saHgVt7M536gXyUalR1Xa9dYLm6TVzd6Z2ClK
J5GpHeAmchj8So3WbyaPmuVYuo3qHiBQ324wXtEpYEMABRLtI6zoa9KJkqLhAJlkkppm/cW5DMxy
+OFh5mzg74bYAcQ6/EwmZA2sro5w+Zlf7+QNtcgOrdDs7HqZHMAhhQxUip5iZhJMIsU61GfQTc+K
wPu4pHKImyNng3rUsfZ7bJN80l7BAs29aoRJscAFrL/O/muS9ro7h5rOLSvxvG8e6Ii0X0IRDuW8
15xEw0CeVtvBx1ZgutbBYONNyYD+YCFm0uRc/Qbp0xd3qgpAhEVZPTh+HL9n3NCfhHQzntRB1SwP
0pLJ1mI8y9GwehIPfhwQ2151lt5bBcZNBRcTibd3E52EMd0gZycL9MXYGrM0wpQXZKlNHCGrZTFs
qktil9BmG1c63PNBsp1/t6ruQLw/estQLq/fuyzP+FUJeMmJCyBNQl7Sr19y+/2vFBrdqg7nFxPr
Ah0uqx6Rkgr8hxPtelIiTqvjz7yJpznXNoYBK0NbHj8NUwafOUeksv8gY1BVEJCWL8sB9RAOl60L
Gi8U7kWkR6OO4u4IYt/wlLeOpgZdsnVPar8voeCMkEWkxqzeR6OQSaxtYacB9N1s1LEjNkzwBLb9
utkeQBnxBfcwAzZ1fmJWGf9err7EkrT8Es44NSCKHwCOanLRrKJQK8FnWvMGrlyooUVSoDz1nW5/
Oyy3kehm2shJYjRw6xB667QvqRIjlbAhYC5BVAaRUMppPCmqIBAQjr/+6v2qenkQiVC2yQ9RL2c0
5XaH0aPtTezgl36goQR84yQO76n271QUI09WvIEirBCTL95fK9iLuM6wvWwX051RnQHtLde8yP4t
71H0LFBMpSbUWbSv8hcJWLnAxKVdM9Y2po/jG6LtlAE2Uz+kuQvL/7gc0KlLlFmNsjAPrKS1j8wM
wysDBKvg6SJoqYj0RajSVTyf/0TQWnfi3/kUYKEXsY39QjNC+hhJ2JZmSCZ146fqZlAKNr1Ybbaz
Xu3VX2HcFB7VF13F3cTa2mwHF65fZWTt4ICog5/L8W/Uxa7gtM/nKhKy7zJvxxXODzpfaXl2cvgH
9KTOg73GkRiEyrD3E6c6urb6etum8wpNu2TcjkSOHlC6y57xjjAH7vtBOrXn66h8nr5KDbxxKUhU
B1ZpPAziS23GX89YjnDRmqjqZkrz6N6PkNkO9eKR3kanBmnd1kDrvMHAZKoly53QgEq4r77MAmZA
Y3nXk80ei22s31+7v3kV4Esiwl8Kbu+PB9RWH4dvwjfGwnhuxaBV5Afj11iYrVNJtQGv6NZZyWvw
3BvAr7PmTky4RSjrB/8ZVTVcShWk/fVh8cTvJkai/gAP541U2dqO//XdUEuGJMFFz5P7r6VdWOPB
90M5Tab6hiHc5rnRg/uwCaP2C6v626nUGVMIQefvMdpRoaZV9j2W6GPhOnOERGzGkGTBq6Xy0WEx
9+SxaMH/p3vDZbs2HaLQcEUyhVxiC9tq5Pngy88fnUrKWkxuNGaqrLuxNGBiqU73zuvlRT0MpoFc
pEH3t33JLcnk6O8MA9xnXyxdgQIJq5FQlMmv6A2mo3623/4ggEIitCnsmhtKy1G/n928CXxRiUwQ
toB00T77BLhJzSLnlvivOIrKF9V/61XIR11/ZlK6u3Kcx0alCU7Co9djtUHezRI1zmZ51yf72oQG
gJ/kQxeM5fGvbE4VLcfVxaDCJjgsUgHkiq03sYJ1l2jkdQkmmWVW8rvehoWyE/uW7Khkb0t2Qr/V
OE1d/JXvhaprmVZXaN1h9whuXc2zIn4zdunb2hnPWzf+clB39SJ3NFPKGJpwMl7gqLciLLfCzavM
t9Y9GpcJXpAnHyjoVi38F/JByqogmnbBsgWPoXl2wI12mO8mxUnyUeIvqpfoWMVXMuKJpfBQOr5i
PfuXLgnuyI/t5KIkJnnEr9dCcme4fwqvkB3+yv3aBbZ/UJBOI+0u5MB1ikExU9qp78HJGSc481xa
W6od49x/UEnm2lgmuWp4US9HAgla6085mHiFNgs5wBX3cGFCIQSUYFAcpE+7tQBWNv51Bn77yrp2
4bK2kYNyzLDphjnslPx3Nv+mbFYP+8mWXxwJJEZEqa/CpVXkhFxeMlpjpi8FndedyKbWuhEUfZMU
BekcWFL7XN17I1wv5odZIox+JAfrIRtu068RHXKx3SxmPkAaLp6LiQjhk852QmDYFOPi1clYGm05
p43k9rdzdJfZWCQGwDxENWtXkMaDUrjBTpPOELJZ/RygZ83W2Y/RgMojfSLr0eNMe3Nc4rDj8tnI
VBh4QH5BKUkg/VoxdzhvaNMOKtH0uqPN2P4pxG0CbpAwdU9sPn+pMGUagGWhBOkmqYZ+jttsn9lJ
DFCzn9rqDknZoYDFI1P0+5rQXluiYWgEnxOXrpPQQ0uDknqjlZ6JZRd9SlH8GJVlPxf1VXLU1cWX
utG/ZZUvAidQofTLcHXxl7cBl5bFPmMq7SgU0081YeG+NZ+3jsPzk36jOFUvpl+aUbRz7ytDUfJS
LLBRX344mvsNbuZCh7nwhcuIs40oGeGTXg5B4Q14De66OpgsXvrvDA6306udBFANVU5Uv85YuafE
80uZTajtvqQZmISNhSJuj060NKA7A4uvw0cHRP73E/6f4+M4iGhaAR1mwUkcIEqWdGbnW9X5Srl0
qgbw9U9uwHq6C4cjzrLLgAcsK2GSs13VGqEv3u+HWBttZvKJ2H1q/4aR0euNWII1SJ3+rFbc+NQT
cWKTwC/wEDXBmz6x68LdYfOUQSdidX0KHls7+i9RxJHw3CaPM7AEMQQmmULkPAomGvf7btMoSDa/
DH5AzuCt9dECYqwR7iGVeFXV68gmTK21WpkbTx61kNn1IOmKcdH57QoVqv9HGjTAvEiE9KzI9/AM
eqRLbTxDNURVZIWkmE0HT6kgy0MhEDBmBhSR/jnzfw/GKlMuJP1z5q/0SH8HOXOl4QtVDZ05nypr
lxxgtO2witdES+qqu4Lxfg+BaQlOyA2NJIP21vkNvppC8bybfNmep57vHtDwJbprJWYpsxMZYK0q
QPpkNodGuXmusOe5WH5KkIidsFwq6FG8gJVGcQdcOBeWffzCL/ieotOkjTOklpjsaB9jktJec08a
v/XVClrMZThNHt5fjfaQym6zF6MK+B63Q8tN5lti/9bYh65Beianf1BC+8dJ/dt3Xpquw+twQiN7
t6oD38hXSwhjqAMvGLGiVBNoUM24tBMEhz9oR9ZROdIbQwy6p0trqXgvde27rOo28OQFe5m3jGyF
83RV/vkiQr69KTJ9yboP4cqUhOa09+oY8GI/uduz2cgLZNpx80NFjoU2w9JW7pPEcC7UovOUsHqF
C+cWuF31PQk8MoEVbiTgXGaay0iVsH/VVVXgkcTKtZM8TAdk422nivqlBDXzxntTToOfNUrGAyly
2iupd2xCu2qFiwFLAqY6SF1octQjvj3nve2U7SqYfws2s7o68cw3wrZGvJTPuc0I3hZLH9TVMF0N
vKnOJK51IlIn7Qf8Wo3u1lUIhiea2+knff9YHBQiFJc/n3LGmnbPNRftRAxU8UtwrfloIa326DIj
wTgoPaiawnjXA2IG9x+cjnmll0xThIvaLt6jAKJ+MSkJywQBW2CLZHGYJFOo1io9vyyy3QRneLfj
iUYmIUMlOTCIKZ/lqd5Wri1ZuMr0jqvDqKVXVGtI9ovx5LhjhEVnD82jP07y4qICMS0gf63/F6GI
pb7wBc8FdPy5WH2Re/gzWLF/K2ugt7+rrEiWTlBkfbQHj3MfjZPPbClCIvoxaAEFGqmulKLcMp2b
A+DLdiym1tEMvH5ew1soNHczkKg6Yf4Rta7YL0clCvrOYkgVzZhuteEbo0sgquvKoGM7/NObaWfR
EaSapO2zzea7hFxPbuBIFkjP9QNBrYfo4Mx5i0KCg3piJnLWXT9UA/lzrkencBC5RyCPVf6/Ng/P
LTESKU0pxuMWsP2UE0odT7YjUEwx5avULikOJYCwxnrEH+hwSmD9iSybUc3aeGf86JTaHaNGEZbq
bgF8BjmhpRC0/Uds8STCyB5TZx6Zrzvclfnd0juB3lj6rC7aKCt4tjuzukDTfrjgH/tAJZeTK7YV
6Piz4EcEZpXDObwyRUEzsvFJgvtpBDNcdzbVLG4POjnLKFTaOWX7LA/K6YAaBjVQQLBRvYvQgdub
Qq8OB2epcKh38VMWDkF7SC7qP9spAzCu6HLd+1MzfOcgMsebckMPG6K4l8w0ps8Ixa6wuL0csSAr
zE2NhysNOd2UsYBHjxBS2gQXCHfewMsyYfF71vYJXZEHTFP/RyLrOPTewkOG9DUCgf43mKGEweWM
7CwuAGdlFQkN8m1+YjdPy9JX7CewodlVecFDzsRgZwjJBcaUBA3KdtLNjxPp5+q6sXHLHRoeszlP
KrEAnystA1H1IKvBul26ko9nA+Sg2qvwd7iKWvYGfjDULzcFWuBFjddPq9qN2xKt2bCpAWshVK/A
G8G+xaAZSbLArVINNCEUgM+fa+IidPwlHEpxwLgQ72vx3nIQka3t33c20VU+ABbo6V0LarnkKPlM
ZCGBtYv1cncAz3+Vp4Od0I139nU9hikq/IvEg9mYDCKWhTQKi78ZPNKe1+XljpTlzQzZ1narN+oX
sLua4PYtd8l1xRzxk5ss9e4Rs1N0Tk3OXW4oB0Pw98PpzyhJMylgdYQdIxKvV0IJMPvtEOq7e5r0
CeeE+Bxg7uz3fiALdLdy2XKBLbUMx7HTcrtIgnQ1k894PW3HQoLDa2VZvgSkZJ8AlRh82lMr/E+j
UNAkkUBbQSYhcxT+VNMYWNUSXv3Ryh29lrHB618VLt4wxKMyHAep3mFR+QdKzufgyCXP+38jNocc
2hAuBt7FxAILHK6OsbE0F9nNEXvP6KanJHTITAoj/9VAzgphWj80QYUe2pcnrwY66PzrKiHUvXIq
yZB6neF72wv/UCbnMB7Blk+0VIhdpIoxwj/KyK+h4HRAFawiqrMKU/CWmVoTC3SZ4A4T3ldWwB+N
JNWwyMdxavdAK6P0QsObq8MV37FwOop0JVZf0h7i8VaYGusxPZFqvlZ/J0v1UKnntYFp1g55jfMl
em+/VQfzv7/O9MXRQGie4DW7tVWulqGlR6U2hntMOXWJ2rHSfMQEdNp4VSmfj5e0heSBh/tggE9K
kzYIrw8RS3LK2hqd1Gk14AGqoQ3740FIN60OVpayeIr85KPlLSI3eoj8vpgjT1QTyrXf7Qy/OmSE
/cxZwbC56iyEbs//ZmossKi0IujeqpytbiP/zQVvtJMDhDNmC0mbIMvSpASz7l6nSVrJ6+SG9MOc
0seO6gCHJHZAjVkaoGgBinOfSpmfIdkrhKIlU1OA+bSmtstBHqatu8orGszRxzpxAukGoqOaJkNg
PTnHy+BwpUvR4QFl/UGvEwOzkirFd56kav0TTKJXF9twPHG8/BRctazu2N5iPJ4PAI+ZyiYqI/v/
X2Cqg9x6XTEN7GUxoIS7xwgvVZlptlWbSRcasl98NIlROfH3PGl2DnEZNC15vgg2+8YnXQXvgFHP
SQ8MWUBA1SKrs3CkR+ROTt2sA1nn7SDLJ1EtVj54Q4s4YCvKw8IrUs+6kK56TAHTtGyiwgZBPQFr
EH6wbaP2OucnZd7AYJyvhhXB2K5Pl2OnVpYTJaY4vvND6/BdyxV5zjCfVHr82gHxwfQoiy6Edp/l
dp9ND7EuxSi8fFamn3JJcf+Iz2ED7F29yzvNlOMqRbafDYkNJAh5LQTrZB57sdvGkdRuJMNkQhxF
tV7B4MvvItvLQ+jhLtCNjZZmR4hvTpQBNvCXVpLy6WIHeMbvf3CX6Z67OGBSzinEnWmBzPsHPh47
nsivJC6YM7czxTfFcvlD6lX665LFJRdc8VPW13YlSWsj1JYQeLbPg+pMVo8Y6+DJJxusoW13sBBG
LmI4hkBBZpFjwqBSy5wkyeI1VjfOXZMUuoFLmHldE0FB0uTLGcHN1nSaBLrursf83Cc1dTpAdFdS
AQfrI+3S820ZmBzugFEqahvCNW9O2i4jGGerzaszTUZ7CXlBwlHIB4bYf8v6li6rbs1K42ndBB1b
XD6qPFAIVG0gLBNhlH8Iihakwr3qosSYDTVIAUIc/xbwsGYZMqalU61BVdb8resySnRViuZNUVox
tXaKsRBsyvfmnaXZBcGxkMWRaaPeE3li4rDswpRzN0YmwGrtllpJG7S3uHZP5Q8WilQdE8WxLfHC
GUf+SVtaWYIECLBNhvms3IpMVgHBMrvEDgumFBnd+7HQZ6lG8S/8Esb2bMJqT6vnKiF4WxbS72KQ
IMGauOLBEpQok2Noy7VdCodUDq3+tFLX40vtr/PWGJGFx0xFqjdqglGHL1KhrIpH75enFjwTv/iC
syvsK8yRZvc8GmJqeNNc4se6RsmdaFz9S/eVn/OI+SnEJVyBiZHOTfL/wNMsfCA0W7OtvBMf1oyy
cYyHLnTCMPj9vB2CIKjorDZk5r16ZGg29QrsuSS1UlOmxQ4Yf8fj4hfldjHWaHy9yw7ub9Tjv6Cc
Lw/GAhx3+mI5gwr5dLGiffKvSdhI9jMjplfYIJ0uboN69odOKFu+M94o/RNmUX+KIQP83sfRJBk0
2qEoYDhiHRLsvZHyjGF4dyLXYm7tWFZINtP/0cVc/Y5NJRfRkFnY9geryAatWvbpn7SoilQawRGh
b6+9Slbrr7ZUZd4VazS9Y1Ik+HwVKJgmi1GFt7hs+GKFP9P4kYRsS6VZRsJ5jR4M7GL2ajd3ObYE
lVI09XAYudKK5jRpfKFJs8D4iEHQ1f0jburMG3Y/osiRcTSeyoJbkKMd4fVL3OcJUv6K4G4DFfPD
1MIJhPFie2pxt2Zsk+wMHt1l7RtcKlYWJhUW5bI8BlJ+ac22/WrLnoE9bqmVPOOCN6DrXoChQD2s
OG7TjZU4OjGVRvQ05mS7XZtk6O57rAObbECF5D85lxX7tdxtfiKNzgh8K+EPJxIXk5SsDFxnaRCC
/6BgiwWebze04xVES2i0/pbKuqsvUigiby/T2zvHJSWtjOx2180Z30t7cawLVL2H+HRqOaZvosvf
eIJa4wfb86St7sPOikAoZVr/FKSekJfCZFJ4bJ5pH7dryDxjONtTliaBZFr5NFMuzs4O1mOFS3dj
6ZWQm2Ou/+7WA9AbPold9xbj9sdu1lPPr1QYhRluOyWU4kjqCaLusbsB/PkqIE0HKUV9cfVRcZwu
a9d1qQsjIFkxOjuOyfD7+t2DvDt2Uj+kEcxjQP1L24OZVZWfn2jTVs7A1AV1XG/glC+Ydgq5m4n7
9TGlBeUmf1uTWHweDMBdMug4L1O6rUOs57sevPpUmr4aAjiURYhS7d3ZooqYvAAbVXcMKz4l9n1R
ibiQ4FlDa5gKXxykbAdjm9hfx6mEfDgZedCPd3RU4nV80nE89AAlOMQVnD8x8yEx9WkUyhifmcWq
6XueYPhlsJA2Bkct/xv74wZ3uTRqmSiWg/RErxfIVX+RTGFTvePjyxsiVlWZeY0WVV5Mwb0ttHk2
mdP5ig0WH4cL0U+RsE5OAMakHWllMWsHec12VwbgZ0DJyaihIN1jXyAKEelzyGygcdCEmEQ159+o
hzu59uimhnCZBBCbCxThyp1CGolW2zAub6zCPKZicnomp+j/vdaluGoaGbeKlgVEm2gkGMjBOQTI
otgB1g0JYzhAEEi5Wox+Bgx6we1Nu512OmfVo1kPfE7xXKyvNJWsT9hXUAeT910DpNr62iw9Dr4F
ARhJXp3sasCgPmDaVJiooxwa4pXvd33ZX/zlwuvaSF/RQdPWrBzIjhd1+9aFU611rjsI4OAhFwuy
NcAL2ys7Q4PFcN1GHEllGsfXxo/ktnlEB837aRKJnyoG2rfjZvjj4oVijLta5F0/nNvkaTSag/5F
y71aa5sfaenXC0gwqUVQhw91pxw+H4/9Bvz/MwkiCg9mS1trr2OEvxQFS4okU/AWm0jTG0/PGgwJ
LT4obs0uDpP8FJ5ybhaf3pR1OWsjcdCmaYLRvIm220/tKaHcAnVV1/N6/gL9uhSrRe3+YqaKAnGC
ZXxL0F0oPoehQonFvfTaSw5AsES/K84E9GJZzZuIXzDvm8ZKIVSNFd9zM8S6MsnjI7B/MzltW/SN
CalaQQuorFijydPJ7FWQen6fNRTvN2Uh3NUq+7KlWaFLz00T1Z3MCVkR3zAmjQtk7Jt6RSYc3bzW
QTr2Z+A7m4B0ZrBI8VxdEru++HVKw+yd3QNjjVkgu4a43X0nc/Kr3jEj4x6gptvTkX9FHZwuMsEd
V4peKT/PaBx++rkMxc3YcqU3J5uoQZ7iAUdlVSeLb598C7WHRpNsN16Ow/S94Q4kB8NyzG7OJbPw
y+RVkb4we7xgwx6/YAXSXcwFo6O08jLDnvdrI/K/H2wddhzTDsw+MNzvb+sOqyYG0YtIC6jpcIAK
iZMxsYUpDhU0uIWVIhveWCtS9BTiVtZ8IwipRDvkPWb285cftH5/3Y03NJQoZvt8d/gPy65gaYxY
Lcfhwi380RbX/YdArXpGuDJuCJeUiUncvmpH0AQezaCGvIvWP1+I1fQaCGUXE22WXNdDnWpNn6D7
F0do38l3G32GC3W5lS0uDU9NajOj/RciLf6zf1I5/o+F8ycSUSugqkzIAuzody4SYanw3pCCzkMa
COdwvUgogMW1p6BKLne/BhR8SKgTYZ2tR7P2ubJbZOwlHwk5FsDPFXMjcApu5GKfFFg30h285IJU
dmBmKGEkvI7Gl53JU1HnP9LupH13zBVn2epaEpEZzCe7+ane3iqhfoyzWjqrmuVsUx4t8RoUYszJ
lNMqAatXzWKaH2NUFDLTG6Ngv8eUwiIap6X4AnOw8LGKRCnhN+i8T1C5C8W92jmce9j7JpDWq4Jt
qkwIOU9o8RtW6KgzPwxbLHE6BmQn8f/5ykqviXJRUKWVD0f0UYDKHpIC8rO5j/gGQD/UOMJ3Jjkt
BpIC0Sle3JffUp0yu5sAWG6XKp5+Q6s8C5MtzK7VjywtRj8OBoifgqrk+msoLFdXUATT5qCEugoG
2eG+tvw+yTegIMb/E1IQ5myLmtuVBa2L6ybLkD38XhI0RAbL2qbb8iDKW1E7u7PVRuMyE5SbRqJa
TfzPL8zBugAJCZEgNhheyEByLoYWcgTloxrjq0V0do4+xdVZIgvpDXodejaBv2EKjScn7EGn64Qx
Rlyd/jZ2Lzg226pfP7Hg9WANWGghCZ6CUbT5iBoUAnk2Dpj1QVZYVhh8C2pByN8h6uu2HeMJ9q5v
eoxc37dg2+XcZzrQCTS2ZlCxQyOo1DTxM2a5CXi5sDz7LDlkJtVBaa4jqDv7Oh4CA6n1jk9azcqE
QqHvtA35oHVFpSctpcV0MzA96XqRSNXfXrBe4l+LXajqdneGtJ3xOFak4Q78YXcORO2tesidY+2B
AQgLanHbg2Qjflebtr11O3jc6Zdsi5zPYxQy0dSto0twajUOCtHum1yYcLIRp1m/sL1Eq3f9ZOn3
jKma6VIqu9NqZXwwif2qa30LCFJHP0U0s+HNVb5NG76FHEiaog4O2kooOK7XDFODM6sVY4Q2ZJLL
prQwwtgOEt53Ti/++BSq9AUlqEtRbAU9GgBI2/CE9IOqLxpusTxltASf40da4cTWfXBDfdQjpu+6
jlBeSi3GwNle7okxt3BHerDTOAQ8Lh5HAZPipV7i5fExiGkz4Uq8KrKazPeamLdvsB7hvIgj3SkQ
70kNI6l2MG9rbn1+1S6WAJrY9ayImJ9fu0uVVpCfe+HbgedntTh/Gd/knLo8yOE2gRnyBpxRq9UW
G6YdScdOxIPU8mJ4h5090Uqv9pJksCs/qddSzl9WXjrUk2zX4ZQVgJKfmVxFzEeQ76gf86FuH0wd
ko2hE9NnWzUHQVyBOKvvHX9oj0JiZ3h8i5MOYJxMuZ1F+TzqgNXBqC7e0e5wmKEMVzyWtLr/3z66
j7SHK0b5RM3/ludB0AeMyiGk/nPr2Kp+hRMHgV60GtekuQ0sSY4ys1MkdOUL2BQNuGSBD2pRTHj2
aDIF2qgQcYqX5OyYiMkrZm6EY1mINi7ZPDS23samnM70YsF234kZYA4JWC87wT/JIRMJh+SbLhgY
HQKl5ccRhDnYB3B4YOpQEkYKpdsLNc4mz+rr0fcRj1gp59USmq4r2Y/9Uf49s0AjJAa80hBqcsMo
HULGsGTlr7YzhR1v8XFVSP/uPQfcszOffl3GDnAXH2vQrLC23BxLig5mZEfZV8RiKc1Am3fVRgxY
T2eJAwGKq26xXcaah9dyiBID5HZufTtxwGC6a6XUfZn4Jn2qQzDx4QJt3UYMbf0aLoa37zG2LBLW
SCymhk7DMG8vPyZh97DxvLJg5bzi7Hecr+l333kFzXFbgxTIahU4DUcfkzmXuBNJquWTEYDlVhTS
knZgDUzcsfiJ/sQX5qWkvj73Qp1XN9M31LoH51QYG652/Gz7GSNwx2nNI2U9ahrg/u5PI1V5O+W8
66dS/uFHVSccd8oY5K8+LOp2zg6V6qjxLm5O3MJ5/DtK69pMVt6FkKRYsJdaTgWf9udymzWHXPXW
SsLjSanWMUFRZ/jhiJmj93K6TN3CylOoSt56GK0S57DYVnBepPhhVgGZAEEppgz6e1RB36PuUFY0
QXorbFemP74A1mgsyQyly8U700IHEIrxfMFaD2dyuCVOZn8jr3OHk/Yuh/AedptAZhfNk5CEefGe
2zfrTY6VqeyJbIPYgy7tPmE5ptnC8+Eo1PF0ymy97/yxVCX60II/P9b/IqS4RoeWmEM5mYpDBS15
vFpfl9qFZ+UDidkGTCMnJWrXUVzlPua9MXJXWykRrxvw9vVLXNPXc/7DbiHvB9f9mfHJuqV8v7ag
BJYEmk3Oi31POq3P4fT8+ONGlC3pOZOUor0g1t9jNxRXGeqiiKr1JMBqstjaiRPEUpz2MGV5fWYK
j13FT7DcAB6VHpjvfNC7GJTtlMFQn41KtO4WAAap+76ILOlbnhJXN8+ic1fEYOTGUhbhkjUSaXNo
kcqKzqaQFfNcdo36tGtP/pVN8vDn9IwI0QCH6Z2m6x17PPtRooSBaG89qaWRsN9TG+UuZmacyVu+
mcR7IsJC9mTaYg3iNB9knGvfnrRyNdg0vUcN0RHVN9HWoQV5BxaO1AG8wVvU891YV7Es6cXgM3xG
cuWw2bVqcYH/g+q5fEEQQFEjzlCbRH2oJ92u7AsGG8LKFpcod9MiKmQnx4ROjwWwBlSMBDQ7AnDn
g9iM5xJfSYTeaZwTKGAw5pfTP+fxDF5ZW6l3N6S3GLImP5FMbL6NkXomdro2SrNNu01IRsZaQWQ4
6DKnvvz115xVGMAoFnWjs3XmFsI/QE+FTAfT74e4Kywj6ClimVNsCLxSvjUzjyzwa//eyuPYoXeg
C1lqiBNO5Kbb0Pq8zN14loyNSdTOupyFZiUo2LPhXYnYW4lOClsTzmBCvxrKaoE7koHYLEbFapnv
HKQ50OB9lDCDTLyShL+nzJ5ciEm63Z5lXCZusKbE5sIb/62Hs05LdoXTmWbK5rDQ3iXF+QGKE12Q
Epee02mnrRMwBQ1r8A2PBwQWIIsgXyu5ELIdipzcNhb7+EyAspxcptwct3guwkyzxWu9NNDcePDT
L6e63qnPdXcrwbo9exc4KNqRVGw15IZgEtnNMDXyLCYAviC9LZZV6A5z+huFsAwfx0s7L++t93Fu
GvQS5gM01jzP/bXV4+XH2Fugssh8rDMozwQsfgXyqSpZ072KZpH3rxwv4xMr+RkLGjBRVyVHEqLd
hmJSYjYHLcf++W5v8/nZZukDLXg7dwlMr6Yyg3ulUOXCoaNbXaXp1zveA+gu8STem/8dLo6GthFw
aIZz+hljGeqOhYqxRahVi2AiZ2F5C095e3G6q3kIzcSAgdtaZVEWS1wpm9YCH3xqqP1kLtA2pnlk
IBfGXmtf1MY+wRmtnsO0qX273HP9YGSUut1uaM5Ts8k6nYXgwykv0+0mj2q3pZV/3dgWk4RiSRrU
CHYu1MH5JXERnfZcyqNb4nRuvQf3UX7sQ39IOpskbL/jX1BhRO01i3srNMGz+Wmr+aTrDjASuV0A
V9jL0xw1fx+5IgYdydA9fpflV5g8yJ+5Vg/hYDWS0xaREEZv8rX1riWXHKIu4QGVkw4UMbTO25XD
DyvHrEX4CaFbjryqFEoW5lHAdUNmAEYPWsSA9dBCTZyaR2V3eZoSQ9feV6m1sGNN5l+awpPgSXYg
64xl/+XkVx2esuQRnEVNGjbP2+5bsl3TiwZCIV/lnZ58E00wHM0LPRfznhnL7cgFV/TzciFXaWRN
wt6yLaqF4E8EZxwsnJ5vUD01Lii3k6ieuGIxwN4px6tmOns/PlB8TE/DXolCc9Es6h8hRTR2uS6F
goPS5K20IGyGGdPly+1ceaAGMsirMlEclCGdEvHpTOoJ5JCx4CKPpAsoPo+R/GyyD0C856qokETY
JUjVna69TxhTaBO/D+YWVL4gZrCwhaH6uqqqWr1MR0C3xWFBCRzE8oZzMBMPK9d4hhu5f/CAnUhW
icZeXFfEJmvJkP3t/uOLYGwi8h2FgvfV9OeqOzmtu6TOt9oOxylNGceH8iyl1raj4YEzDQIYtMol
TTZsULv9C8sE8la1GG3o8ZKkvyY/yIdsCEFGH1u1HM9/40zOJGaqTv6XqI9w34jhO7cfpvaVQV4n
IfMFKxc1h/bPzWvEldmq5s1JOqW31d4/jYWMGV6pJ2DToWlVxXr4Q6c7P/NT5yy0mS5fuGMGGI+7
cwzF3bVt0hKMLLIUVv2VgkQeYi9GH6+YQ2xRmLdHV6R1hHbK8Xl8PDoUT3NNwEVrBcXCvXJRg9G3
0HpGIaCDICax422dylEuInIK0ELBkku9CJSIiWz8dYtJCXCeWYNVKkE0DKNWqxKYf1P6JcOqxvF2
HcAYAKQOv2m+fzdbdxpQhyGTx0bEyrWCCLzdYBOu9Llw20gAUPQPEmRmn8TJ7ImGQW5XTf8e7aHf
ylKqPc1zTseoQiBrxppYMQdoDBjKKeLhfe9rDyRkzDthDNZfmH8LQZrkJt7YxnowfwKUhr6h74ka
YPiFe5evonRWmna6NteLw020CdAUAHU9U7k70crYP4/1+OKh9hotCghJhoSpWyNJVtgXAZY3zkQB
LIpkAJ/cd/ZWohr95B8D1wiJYBNVm2fJ5cAKYHGWecGUxNjhIZBQQQ6PRE0eOIOl4C8qAPoeg+L1
w1QOwARZUTwtaIDDw+mX+RLBpE+n3IB+hshtFgprTd5T0DRgrJZTllnWHBjPnDWVxnvGb7A/FzCx
+xxWx8mNNTuxzwkDledot9aQVbW2LdZ4YV8PnzNr9V9byRSzJ2ADp75sUHtmDrgb6H3sH/FDwy8/
FkHMTCxDq6b6wldRjvvq4mnlNAfpIe/bY2V9rDxn7vVXB7Z0FjNXheB29stnUpCM/WiVvAq7+Jr9
CTqIwmd8Oz+nvBsfDVpGCU5yZJOtLGoe60W782V1MQmeLk5OtTw3uVTADwsF4RgvOlIvrslzsWMC
PbqXEpNOyxSfes97l7kotePUGspOH8lwyvESN95KKr4AV1GyDSHSlzEUqGDhUvyYqQEN6CV9sNIW
z/pDudpCBLCtoAoS+c9zCN0mL59vpRJkahJV+czshC3c3DLTxoJdiShUyQXWxB5WBWMipvW4WbsC
XqW23un2Rn8UDc2Oq1MLAJwLHAC2v1RBS79W78bk7Iy32Hn6bVjhlZG5orkSqxh3Bjctqusn3or0
gcm2hmEZG10ZLqnxdyC6GTykg3C+ivF1KC7sF4iPUaAuydZ2Nx1SBNOvFBUoagbAfpTPn8D5tBRk
1EjdA9z3o75p+UMZ6J9G7fTp3N2pKmr0dcIVsrQT6vtAWIN8LT5RldkaPJILr0hVdRAtmBdjSU70
DYhBaO8jINMrGE8lYmXqsuFVYh5LBHvFiA3qolzG2tT9pNcFOBJsS5i8PKuW0Fxtk+Zd4mkWqXi+
LmSKrjPuxGqHTmyFGEdz469hG4pCv1U+CxqE+pXR+aORyXmhE66PzhNDhKONT/eujIt0IoN1APhM
yyK4cy2jZdm/ok7KtqKQyYMRsaH40pI4tlK7cUZCrBbb6sZgj/0SKfmZAGPO39bE6jR1mEYIAVm0
puvfHbQh7oio5pmNbq0gULgosQH+Kkp3YFe7Q9emxCQVln4lpIu3lCnIFgogk/YxgAnKjkes98gU
bZ71iGfXa8u5ZTA34TodmHHlYju9mCJY85WRqADepu11qIjwBYPKlMuObgjZT6SOHZtYAhmzmt2d
F8jQdKKmMgkmq2WQDJW7+sP8uF+3WK6+MpnY5CuscIKlt1NwHz5xKbJFziM5GqFWyQ9luPZbMDzA
lW8Mly9MZJK7vR2w0j4iqLRBIcCj3XP0yw9H0XoE7hTsEIzT0vDWQlE7ay9XOhoSZ2N3d0lXeliE
LXXaK0SXR2KvI9vaoUVck+F7bOXMTKL2Un2YVVDEJNf45s8ePE0886Qdv5uEiEIVOO0PVAUkIr3A
7DeMtbEoUgSrnZv7a3GD4otsIGAs1yPF45CGsWfYYz9ICjtYPwCrQW7f3AF5iExTLLPE7Qj4Qv2l
TH07AfYQpqYi2fGcodKL84iWXV/0gZ8kAPkQabV4grANNMGnXWd44dgLAQo34NIO3uAZdsFQvHCL
lK6BZCountUE6T+FK+TsbCBKGZJgmc86Tjw3RmF4QxcBtJH6MvzatsVWOEYWZYuRbn7fY7YCfO70
66oPNsdTBX1NKyKTvm79hZgNkG1mQ9QHa3Zq327rcqNhtvBxVrgoIAXtCWOmaasaTQG4rTDBWAHj
8Olb7duYz0gbUSHUQupXmsg2gG2hfqN+47hi9JPewmrMaY2O8qV5LJpKzlxqRTQBgB4IlCTVQaro
d5gFKaOeCHswvmlmRQC6FcM/AUFRBqdRMdfo0AMbTdlzcCOsXjJSIq/OVv92vsi5DPaIOU5qhxKw
+BM07p5q0HTw1r2ORC9qCfhz5ontTJtWGBTKkJ5ZX5b1/aXbzcKHZDnrJyRNhs/SWIOVfroVr2hb
sDejaemFpT/fOA3x1W0QWKRXtHZk2r5OqijgYDPFNDmqTJT7XYzf2ZykPEOJ/VcyUCDAKvN7DYYT
y4mecAbGLuuuLdmwQjTKFSU5fNGeQ+7/pveIGSVKBp63eRQEfT6b3mwrXkXE9SRvkk4LN/gMShTx
e3L6JM5UXR490JKmF24CX7WPqPDx9Jtqt7sjOSBLNMP0WZ9Ukr/+pIh291BwYzGoWgPea4lLJ5by
byRCHE9YwMVabV3lFHFyeKIe2NGnRIgWx5wE/fV03T/xVpm2wIkit84Zg8gTazYB38vanNmELKHq
HSCgdV9sTQamafNDuIkN2rUXerDvHDZW8KQ2QFzPi04vYYmUAB3HGMN9h/9CaZ/dQ9goryFL8Mbc
cuuoVAN11/02m/axw3tsOPuHMNxrJ7nZ7GYM1lRiTU9flIUvLuXrdwHVZmV+0gZgVNv+A8WPYTZs
PcmzB8pDezk8G+HMrzVZQW0MSN0LWolKXqMSAk0MU9+8rq2dSvNN/4mmkUF0ke6uU2r6L7VlcW2g
cAbOPf290w3E6MGsVXRVrdEk2OO4kIB5hv98RYMS81f8bv0TllCqL1VNn8QQp4pJ/t53zegCKkjz
DmoAA0ZCmZ898Y1P7g/ryZXLytGInfVHgemKy/0BEh39EM3PPIwCaIgWqL803M3tcbh9m9vHhJ4L
NQKHB9ePpqm2lpN0DV5GD5SrjsE7D4Li21UyrwVmTjwTe37nDh9vWTpNRYtDFIMcf5asjwtfQoXU
1t8h4MJAJpGq/OuwJ7AEWMmOZVcEgygZTMTl8+cut0k+N09KbNM3xog4ebgDtc8tXWPFY6zAjhpr
8g4PoMniI2HT+6mJgtz2UUDiJPuPUVcYIdLr96g9G1RzaSvKV340G9MvYmgp+XYBQopj8EBS+K8p
3MeWCbN6NWyLuxlxvOEl9M2xZAaVOa7oWrUVQvdyjulEOVLKCE6V1+4AcnsLT75aMwbNFD1J6dlF
mbEbVMKO4C1Z0OI31z6TdabbQ7lXzLigc6HpEslVUbEMujBVapjId2XT/Ompb4Ya67T3eP9D26c6
JowaTK6MnprcDHBXp3vdHz8qS5s9Ws2sZzBoxm7nMMaW9Q40+IJ/QdV1Ms1mpwzSOXnlhKwNiR8G
k3NorYmZvgAtlMcCHvcuOPE326X8dMKZRfcZXAawEuzdrsQzqFGE4r32rpzWPnSmxOmcnNCMHGW/
UrZLJAo1AkDfOMIKiuPu5/9ocOZRZS8WJbNzDeWujfoKwjJOVHuAc1lpQnCvmvuNhhIbGx+RHILK
FsQgHB1p3UbqrTiVyDrIQB79VgiAiOI9gCHqymzUSzNUqqli0KaOLyWf5cD9VMPtICy4xSiBIjgJ
fRztYdpa7IIb/SRvvb4I0hoVHZmg97HUsIOrC9xV6BsJ4j3gw0rlshokILBXy3A6xyVtyTnDHi4s
8Vxcv/iaHJ2GMarU+v3qdpSqjNHLGXnhxBnypT5l3WKJaorl/+/QKTSirDeJRaaOtMKg04h8isWd
jPgSNpCCV4GXT5YieN7Dehrw0yWN1Tlkv27qeZT2x9L+MrgsHheXBIq+WJEcSaNAcU0qZO0ZWqBG
OrAJSO+niYCzzlt+tJiNqtImtp/LfYvhk4vOa/qrOKRjuicRrkH8A1EvsELAKHFdg4i9eXxel7mv
su0DJe2pFtOiHvPP3gDOo3UjCTd2Trhh9RPVyLypLRTAmGQSsiCdwopFTNhlycAGaeeJiMb85Nhi
Vng65JKeJgiuNUQm2Xsp/2UZHX+wOc+j8AMmKyOdbSDdzV8xx1YIoZ51iYhtNGjMZ1I/+cI/e+Te
Y4lGeNuWCR9Tng1bxP5W3pVlXpF5ibB581v2HhgFKsRipwzIwgbWXfDz1ezfQsxoekwCAMdvYp94
p/XFOSE2FyeJWw6kjEXv6FM1IPi9PICKb+Cv0Bn+ImPlcP35eyR2b8FSp78QhHmGUyDsmI1556eK
6L3FpxhjDIKydqDTyg/lA6KkMPp4sXWwNW+PC+ctjpszFBNKL4phmU6k5Q4ALVGoNDC3Gvei0wBq
XCtFWkMCUtBEHIPIDsZHJGCerPUWkqYQcXFRouYpyV3qOaAh9WSSkr2NqoJPtlEfeodM67z9E8FC
G2CSX/W3oyb3/qXzftyLT8G3LAgLFtHUScQHaeTzyzAXQj3XXVNSwAYlfZBedcHmw32q6GOUcwWI
6MHFYDgYg+iyzCWYIiBsWoJtcqg6KSwCI820IMg9ExirNG2PIE3UaTB1Znlh7ET9R/VBtImaBMCN
8fiX7+E5XRGapKzkFSk/z3O8x6XhNL7IZsp5ygN3kcfyx4IgB36YnZ7WeHPtiUepwPnIGqGPsqC8
adi92Eu4gB/sXb8vYQTIa6yvPym3VRzj+xC3i4u1HNyugcqYISCQXe59yMi+ahmuV/UDuyG41ryZ
JazaZAZ52nzZtOAbSM6mTDvl4AaR7ubRcyWgNW8HWhIjK7Ti2YV949721i4RILbK7gmR8L6zJGBF
s27CgcwP05CDqagTehT9iXeVFrQpi0HuG2K0dKoaaX1D7IlDX2drqtSKb4vnl64NrVviNRgxsg6j
bdlQFTee1RRGcH8/9m0yQ3Q127RaBs5fFgC1WjvHpMMrlrvc2UMeBDHwfSncjiWvcNuAaB6Qkoaa
9N8D4hehm4xJzQLY6E1zlZDngzkN0W5fYK8kvRd+oIPxkVLz5r1t7QJZK9ytobrdVP10sVN9X1Bh
3eOr4pbPAjI2kTJI+g3lAKDR0xcfO079dS/QATsw/kuUOQj7DzrA/bU4FWXD4szUnqz6NIs36XcF
oCJvqbifzQLoly2QEU5jztk0j42u2UMK2D0uN4b4wFrnj1/Y1MYz8Ft06oDpWB/g8HGDzbh03oO7
I8KVhNKnfnlqRMQXF18Sw65i3BsdQse5/YJRwixdReb2VeDw4aoYizxwB9hCgdtcYHDvyhyIk/7y
3gi1wp/FKGJhksG9Sx5wa/oMKce/JA/rJq9hTp4MGZmjNRKu+89VVDSfF6QSzOxtGE6zoqNG8+o5
cN5e+gokpFL15ejDN9vKmOs6wRt5zlWfkrYk38FLeWAmZ+WKrguCy6pF8MG7x0il3pmmaKbew9zI
BmqVXyeQO6jQOoEQPU4s4aT1hqfhvF8JCAPi/TDSzsj9o/4hC/tqWimlu0Fv4r/gaxHxgA6d+y07
HfK7XzNFMJ+TMtXKeEtHsvPDrgw4VxMkbb5+mg+vmCITG0bDYP8wnW+1vnkcUJjhhV7fmgX7JExl
3U6pQB3RAtPS0jOntdaOxssKo3NothUgIYMZKXRzpZ29HZbqX9kFLUN2GArAj28rNHSTEdowWTq4
urygdbV0j/PdmYy825vJ6YLLiQ+EhQoeIcJ92JWNhngbLi13c7M+TRRA4abSZcdnAJKxb2AmDy3S
bYv21pNW9mRnjwTp6enmgIyXIwkDtN7rp/Kl6iBb+lfWCWzX44A0gHDJSkIcEaXOSbHpPBTiGdFK
8Aki/q/Fg4YjDUMsGUhoaFKiVMFq0cwDY/lgvaW9wYUWzgiTFUhGFDSd1OHkA/I7bZX0gyLr3oRE
FG9MQb/BAlrXumg9KrqyuobFYck24jYcwmV81GQoYmCQL0yKVRejd6REfBPn0mAQUbIWXlJ5HiNy
+r/X6u7Pehwov//keY6f7YIcSlHHCWjQcx880aJClcqE/fwGY2Hvnkpqpgys7qs2HXknHWIKwmxj
GZo4MG67WUcwQ7wseSG+d2OJ1lWUVYdhVdAvDx2BLgjs/webeLWJ8g8lNJKH6GrkeTvQyS64OBDQ
Drqu2NUCu7J/47bLtBQlbGvP+cq8yyf/SSft3K04bc1fExdCHmo/rxHBCpBhPOswBym94lSjfjE+
gy22eqRiO/NAg+nG+CvP4BpRv0dRSAqIyinDl5yjA/SwbmUFdBOZMzowYBaLiRWmhOta2p214oqj
5pzjUNw2SPVdlAxhxpEcwZcSdi/gz+qsH4ad1QxfMM8iqxsW2gNhiy5YPqlb0s1Vtws6Chkb8aHk
/L4gdYXWesSobV9955pY6eObbCF1xE73NvpDDk0oX8I+5nNTArQWP4s5DnzUZQhprkisfQ1vhObp
DphJYIlXq1+ldnv9uk0G4pVcCNif712gqufNl9H3240ozaf7nh+CBsgctz13djVy1WhadhSQf/UC
2S24OjeWcwbgweKFixmwUoKvwyhpw8DYClfuhRrfeGF+dwR/80soK7KLHC1CLg4tsUL74226qY+H
CEZ50RcPVmOLlE/w0nzfMZGY0EY/PDVaOquK4ZcYTeGB9hMyViqTiYZh4b3wafVtAlRaGAc6JIok
sb3sbcjo5tHXr6XEP74zsIKrKIskP0yLL2AQNZOHbYMWf3OWaSv2ic2+Lu67j2E5+NCvtDT7us7o
R8KEGToUlrycQOJ0lWH63Cqd9E6bPsmtWdNP57jEPrw9Ufm+P0GRl5cUsKg2P7T9bVOvOAprX8Fi
tXcbv6hWA0z8EkeRtKgEl6EFO5PWnqITFIIO62Sh2NwqtyGTLCRurmrQ6ztHc2QfP7T4VtZddQW4
vtQ8M/ano6BZCt4P2WMo3NWLyZ367wSTMrRO06znUeBsW6ZotQSw6ZmXFl3wnpMy/1HJ0LyidhKt
itM7arM05pex1gg7UFUP0CwdCIuVDM/rkFBSuqFPxmQh70yZuvc1Jmj8WQHZfLeX1Zdj/E6kj1wq
cZx0zpJqaZ0k755q7cZ2FyBOZKSqsPxUpsdPSC+xYwc/I4763KRoFeVYcJDVk5gT3eB+seDPogML
Vkvkm8IEMk9bukySBl/gY5guec9DTLoKhmixqA2XZClCrpLHVIQ9eoL/tnfwZBYn70agLXd/FjKZ
IDQJkJ4lwg7WbV5sGJn4pQtbhzU148LV/DxAOnyn70qSBiAIhYCiYwwx8NP9+cQfe9fnucM9e6se
DgJEIWhULLDa1KKibUyPvpjQUj2HkVcURsoIG5Qx7wDVumh/gHB2zzBAJ1sJYT+F5KRmo3xzmu6e
rbThOVnvzs0fBA1UnrUbyAUmPnAtbQs6VlNGYCsULguaTuI0wxxFbhpUrthpNVYCoE2YzkbQL9dP
SVMwq70v9k+CUOPecp56LnlAUBvSqfhGQjsiReuVm7JIyG9Lq6FyGSspCKzJ+g+s2u2d+E8QHYqQ
57/F8QVOrXHwcNH78N2I7nm8/ePCdDKBc33Zb3LJ05l0iP9NLhsSxCCO4jJFgqtwc4SBv+DZAymy
5J5ckBkgaJI3xnUfqLlPchZHfsRj1xFXUhe2nQdI3DEgFQLocw5c1geD4KNJ6eBd9LshPmbGmEHG
fLRS50jP/wT4L1B755at/3lokyRPLctzcmMaIaGjDq3dhwmTtCRGXmJLleKJr4eopyAcCBMnetXo
no3iWtvF409b6xvcwWff9eNJxNdrSueeVtRaGmxtJtV7vUQzKhWaMsAevDil/2RA/VP8Qde5rEZU
ovqNl7Hikp5gkq1HLiSVtyQenjzfKwmCluilwxchSy6VMcqAWMO+H8qYgBHcXTidZVUG6MlGdwbJ
ZJTY01aCQlP+GTzUIk3tV4audiHv5poRS/ivStWCuC7w8fkdFkYClSgwp7COaSM/PwEEjpM46wQr
tahOo/yw6NXOELCLNABmF8jEfzVZwAp9DGRIvrtwQGOTRBdaXvP4q2/98QW+8iRnXmfc0SLgVtXS
aS43ifjd0UmQAB/B356X9q6c5VqjAsAawhgoD6xpnX3u/dxPr6HTmnx1H+64F2BpIpOdfb4xQSoU
RpLCyF9XD69XNmKp/JDF0Ws5Ey4cWdM8N8F4MScJqlsYy/X4jdp90BP6DxBy3VLptcqviAXxhk/x
pIKaegMMwvvoPbvY7kVNNa/NV0vV1p4z6S5qRvz6ElHtbj93SaQAis3aSKoqB3SvOq6Exkc18cxM
PFKuY77MYOBLlz6RivQ3rpEppQ5HSCaawf0HmGEmChVqTilYJ7Fkb8qTPwPrNlWKxiqNysSXE+IH
ZfZGxWL1Sj/eOyZYZ4NQVc3YKrJS1gB1H2Fap+rAK3fwtQgkEh/8jKSI/VBXfV4g2ZXpXoEdQhWM
TpLRbRGyfvryJcahuMe1sQCGus9lCIRmn+71053NbTjXIm1BT8uOQGe/KsD4vckEU8/qMSt7GkBz
PmZcq8llDwBclLdvI6VGmIQ78KOj+Mn1nsZgt4UvT62keB1BQ6bYvxmG3gOgOoC7NA0zjoRyVzX4
2mD8XNaGsYIEB6Eb9SfIJEfSmpE+ICOAbzaMBlxhw+IfYmHP8Tb80X22/18u7J4uVPV7D2l+tqAy
mF0mx8bPAY+QUDDP1GFvIFI0Jrsd896FaCwNHcxlZzUR1MVP5hRhJ3D1w8tkuPE3RifoYi4r+Bwn
/vsvUGYq/Sn3io7ANZ0X3N3115E+l7zQA68VdAB8fD7PZgRv89NlzdxrLvp4qq2yhWrr7vShK8zY
sOLiCYymz/lX3o7RDHzu7HRKfjTwo0u+/DndFumKiYFdkf1OJ4uoZSOuh6VXOqyrWDgeE1/cxtzC
ClEqIAKuRir0dbC8P+aUKWZNCqUvNBMPlFJ+IZ0BqaX17WkFNphmdRre0WzApdX5tHc+gIrT0wT3
g+X2KeSWcrfqTwRp5zCUFzDZ6Ct6EeXfc7Mg2EjBaMeSxq22nKK1PoPfN/PmKzl5PxsN0cL/FglU
gifjrDvrYkEnfzkUyL9PE+fB6psHUzVY0oEzqyidq5L2fEXuac+ZEhnlUH0AwBCA5LoAW3shpct6
vRii4GlyngQOgCVF1OAqJOu+m7rO1qrphTfypgrvrU1oD37UvlFzoSIPBIf10G0Dc+BDCyjVJWAx
R+yIvI7QWN5YAB1LbmYlUsZ6s4TUrt8fymhm74g1U9t1+NXmgpVuL4HswKee3Gz0RyMpaldW7eld
RDZznN/sz2wy0ktvwK0LNLcOKhBL0r2j0iaEWmWpq2l5oT1hCRXcSjNknkIxu7P54snfsw09AK9L
mHxXVVDA6XjwB3cz7PKHQSdXqttUHgRnctDfsv/Yzfyp5HohxOzXu+1RfEWFajzDdyZqKX3p/lkG
A+Z40VRyJjsIsxaH
`protect end_protected
